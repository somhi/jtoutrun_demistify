library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"ec00001f",
     1 => x"f100001f",
     2 => x"1e00001f",
     3 => x"c848d0ff",
     4 => x"487178c9",
     5 => x"7808d4ff",
     6 => x"711e4f26",
     7 => x"87eb494a",
     8 => x"c848d0ff",
     9 => x"1e4f2678",
    10 => x"4b711e73",
    11 => x"bfe4f7c2",
    12 => x"c287c302",
    13 => x"d0ff87eb",
    14 => x"78c9c848",
    15 => x"e0c04973",
    16 => x"48d4ffb1",
    17 => x"f7c27871",
    18 => x"78c048d8",
    19 => x"c50266c8",
    20 => x"49ffc387",
    21 => x"49c087c2",
    22 => x"59e0f7c2",
    23 => x"c60266cc",
    24 => x"d5d5c587",
    25 => x"cf87c44a",
    26 => x"c24affff",
    27 => x"c25ae4f7",
    28 => x"c148e4f7",
    29 => x"2687c478",
    30 => x"264c264d",
    31 => x"0e4f264b",
    32 => x"5d5c5b5e",
    33 => x"c24a710e",
    34 => x"4cbfe0f7",
    35 => x"cb029a72",
    36 => x"91c84987",
    37 => x"4bddc0c2",
    38 => x"87c48371",
    39 => x"4bddc4c2",
    40 => x"49134dc0",
    41 => x"f7c29974",
    42 => x"ffb9bfdc",
    43 => x"787148d4",
    44 => x"852cb7c1",
    45 => x"04adb7c8",
    46 => x"f7c287e8",
    47 => x"c848bfd8",
    48 => x"dcf7c280",
    49 => x"87effe58",
    50 => x"711e731e",
    51 => x"9a4a134b",
    52 => x"7287cb02",
    53 => x"87e7fe49",
    54 => x"059a4a13",
    55 => x"dafe87f5",
    56 => x"f7c21e87",
    57 => x"c249bfd8",
    58 => x"c148d8f7",
    59 => x"c0c478a1",
    60 => x"db03a9b7",
    61 => x"48d4ff87",
    62 => x"bfdcf7c2",
    63 => x"d8f7c278",
    64 => x"f7c249bf",
    65 => x"a1c148d8",
    66 => x"b7c0c478",
    67 => x"87e504a9",
    68 => x"c848d0ff",
    69 => x"e4f7c278",
    70 => x"2678c048",
    71 => x"0000004f",
    72 => x"00000000",
    73 => x"00000000",
    74 => x"00005f5f",
    75 => x"03030000",
    76 => x"00030300",
    77 => x"7f7f1400",
    78 => x"147f7f14",
    79 => x"2e240000",
    80 => x"123a6b6b",
    81 => x"366a4c00",
    82 => x"32566c18",
    83 => x"4f7e3000",
    84 => x"683a7759",
    85 => x"04000040",
    86 => x"00000307",
    87 => x"1c000000",
    88 => x"0041633e",
    89 => x"41000000",
    90 => x"001c3e63",
    91 => x"3e2a0800",
    92 => x"2a3e1c1c",
    93 => x"08080008",
    94 => x"08083e3e",
    95 => x"80000000",
    96 => x"000060e0",
    97 => x"08080000",
    98 => x"08080808",
    99 => x"00000000",
   100 => x"00006060",
   101 => x"30604000",
   102 => x"03060c18",
   103 => x"7f3e0001",
   104 => x"3e7f4d59",
   105 => x"06040000",
   106 => x"00007f7f",
   107 => x"63420000",
   108 => x"464f5971",
   109 => x"63220000",
   110 => x"367f4949",
   111 => x"161c1800",
   112 => x"107f7f13",
   113 => x"67270000",
   114 => x"397d4545",
   115 => x"7e3c0000",
   116 => x"3079494b",
   117 => x"01010000",
   118 => x"070f7971",
   119 => x"7f360000",
   120 => x"367f4949",
   121 => x"4f060000",
   122 => x"1e3f6949",
   123 => x"00000000",
   124 => x"00006666",
   125 => x"80000000",
   126 => x"000066e6",
   127 => x"08080000",
   128 => x"22221414",
   129 => x"14140000",
   130 => x"14141414",
   131 => x"22220000",
   132 => x"08081414",
   133 => x"03020000",
   134 => x"060f5951",
   135 => x"417f3e00",
   136 => x"1e1f555d",
   137 => x"7f7e0000",
   138 => x"7e7f0909",
   139 => x"7f7f0000",
   140 => x"367f4949",
   141 => x"3e1c0000",
   142 => x"41414163",
   143 => x"7f7f0000",
   144 => x"1c3e6341",
   145 => x"7f7f0000",
   146 => x"41414949",
   147 => x"7f7f0000",
   148 => x"01010909",
   149 => x"7f3e0000",
   150 => x"7a7b4941",
   151 => x"7f7f0000",
   152 => x"7f7f0808",
   153 => x"41000000",
   154 => x"00417f7f",
   155 => x"60200000",
   156 => x"3f7f4040",
   157 => x"087f7f00",
   158 => x"4163361c",
   159 => x"7f7f0000",
   160 => x"40404040",
   161 => x"067f7f00",
   162 => x"7f7f060c",
   163 => x"067f7f00",
   164 => x"7f7f180c",
   165 => x"7f3e0000",
   166 => x"3e7f4141",
   167 => x"7f7f0000",
   168 => x"060f0909",
   169 => x"417f3e00",
   170 => x"407e7f61",
   171 => x"7f7f0000",
   172 => x"667f1909",
   173 => x"6f260000",
   174 => x"327b594d",
   175 => x"01010000",
   176 => x"01017f7f",
   177 => x"7f3f0000",
   178 => x"3f7f4040",
   179 => x"3f0f0000",
   180 => x"0f3f7070",
   181 => x"307f7f00",
   182 => x"7f7f3018",
   183 => x"36634100",
   184 => x"63361c1c",
   185 => x"06030141",
   186 => x"03067c7c",
   187 => x"59716101",
   188 => x"4143474d",
   189 => x"7f000000",
   190 => x"0041417f",
   191 => x"06030100",
   192 => x"6030180c",
   193 => x"41000040",
   194 => x"007f7f41",
   195 => x"060c0800",
   196 => x"080c0603",
   197 => x"80808000",
   198 => x"80808080",
   199 => x"00000000",
   200 => x"00040703",
   201 => x"74200000",
   202 => x"787c5454",
   203 => x"7f7f0000",
   204 => x"387c4444",
   205 => x"7c380000",
   206 => x"00444444",
   207 => x"7c380000",
   208 => x"7f7f4444",
   209 => x"7c380000",
   210 => x"185c5454",
   211 => x"7e040000",
   212 => x"0005057f",
   213 => x"bc180000",
   214 => x"7cfca4a4",
   215 => x"7f7f0000",
   216 => x"787c0404",
   217 => x"00000000",
   218 => x"00407d3d",
   219 => x"80800000",
   220 => x"007dfd80",
   221 => x"7f7f0000",
   222 => x"446c3810",
   223 => x"00000000",
   224 => x"00407f3f",
   225 => x"0c7c7c00",
   226 => x"787c0c18",
   227 => x"7c7c0000",
   228 => x"787c0404",
   229 => x"7c380000",
   230 => x"387c4444",
   231 => x"fcfc0000",
   232 => x"183c2424",
   233 => x"3c180000",
   234 => x"fcfc2424",
   235 => x"7c7c0000",
   236 => x"080c0404",
   237 => x"5c480000",
   238 => x"20745454",
   239 => x"3f040000",
   240 => x"0044447f",
   241 => x"7c3c0000",
   242 => x"7c7c4040",
   243 => x"3c1c0000",
   244 => x"1c3c6060",
   245 => x"607c3c00",
   246 => x"3c7c6030",
   247 => x"386c4400",
   248 => x"446c3810",
   249 => x"bc1c0000",
   250 => x"1c3c60e0",
   251 => x"64440000",
   252 => x"444c5c74",
   253 => x"08080000",
   254 => x"4141773e",
   255 => x"00000000",
   256 => x"00007f7f",
   257 => x"41410000",
   258 => x"08083e77",
   259 => x"01010200",
   260 => x"01020203",
   261 => x"7f7f7f00",
   262 => x"7f7f7f7f",
   263 => x"1c080800",
   264 => x"7f3e3e1c",
   265 => x"3e7f7f7f",
   266 => x"081c1c3e",
   267 => x"18100008",
   268 => x"10187c7c",
   269 => x"30100000",
   270 => x"10307c7c",
   271 => x"60301000",
   272 => x"061e7860",
   273 => x"3c664200",
   274 => x"42663c18",
   275 => x"6a387800",
   276 => x"386cc6c2",
   277 => x"00006000",
   278 => x"60000060",
   279 => x"5b5e0e00",
   280 => x"1e0e5d5c",
   281 => x"f7c24c71",
   282 => x"c04dbff5",
   283 => x"741ec04b",
   284 => x"87c702ab",
   285 => x"c048a6c4",
   286 => x"c487c578",
   287 => x"78c148a6",
   288 => x"731e66c4",
   289 => x"87dfee49",
   290 => x"e0c086c8",
   291 => x"87efef49",
   292 => x"6a4aa5c4",
   293 => x"87f0f049",
   294 => x"cb87c6f1",
   295 => x"c883c185",
   296 => x"ff04abb7",
   297 => x"262687c7",
   298 => x"264c264d",
   299 => x"1e4f264b",
   300 => x"f7c24a71",
   301 => x"f7c25af9",
   302 => x"78c748f9",
   303 => x"87ddfe49",
   304 => x"731e4f26",
   305 => x"c04a711e",
   306 => x"d303aab7",
   307 => x"e2e0c287",
   308 => x"87c405bf",
   309 => x"87c24bc1",
   310 => x"e0c24bc0",
   311 => x"87c45be6",
   312 => x"5ae6e0c2",
   313 => x"bfe2e0c2",
   314 => x"c19ac14a",
   315 => x"ec49a2c0",
   316 => x"48fc87e8",
   317 => x"bfe2e0c2",
   318 => x"87effe78",
   319 => x"c44a711e",
   320 => x"49721e66",
   321 => x"87e9dfff",
   322 => x"1e4f2626",
   323 => x"bfe2e0c2",
   324 => x"d9dcff49",
   325 => x"edf7c287",
   326 => x"78bfe848",
   327 => x"48e9f7c2",
   328 => x"c278bfec",
   329 => x"4abfedf7",
   330 => x"99ffc349",
   331 => x"722ab7c8",
   332 => x"c2b07148",
   333 => x"2658f5f7",
   334 => x"5b5e0e4f",
   335 => x"710e5d5c",
   336 => x"87c7ff4b",
   337 => x"48e8f7c2",
   338 => x"497350c0",
   339 => x"87fedbff",
   340 => x"c24c4970",
   341 => x"49eecb9c",
   342 => x"7087cfcb",
   343 => x"f7c24d49",
   344 => x"05bf97e8",
   345 => x"d087e4c1",
   346 => x"f7c24966",
   347 => x"0599bff1",
   348 => x"66d487d7",
   349 => x"e9f7c249",
   350 => x"cc0599bf",
   351 => x"ff497387",
   352 => x"7087cbdb",
   353 => x"c2c10298",
   354 => x"fd4cc187",
   355 => x"497587fd",
   356 => x"7087e3ca",
   357 => x"87c60298",
   358 => x"48e8f7c2",
   359 => x"f7c250c1",
   360 => x"05bf97e8",
   361 => x"c287e4c0",
   362 => x"49bff1f7",
   363 => x"059966d0",
   364 => x"c287d6ff",
   365 => x"49bfe9f7",
   366 => x"059966d4",
   367 => x"7387caff",
   368 => x"c9daff49",
   369 => x"05987087",
   370 => x"7487fefe",
   371 => x"87d7fb48",
   372 => x"5c5b5e0e",
   373 => x"86f40e5d",
   374 => x"ec4c4dc0",
   375 => x"a6c47ebf",
   376 => x"f5f7c248",
   377 => x"1ec178bf",
   378 => x"49c71ec0",
   379 => x"c887cafd",
   380 => x"02987086",
   381 => x"49ff87ce",
   382 => x"c187c7fb",
   383 => x"d9ff49da",
   384 => x"4dc187cc",
   385 => x"97e8f7c2",
   386 => x"87c302bf",
   387 => x"c287c0c9",
   388 => x"4bbfedf7",
   389 => x"bfe2e0c2",
   390 => x"87ebc005",
   391 => x"ff49fdc3",
   392 => x"c387ebd8",
   393 => x"d8ff49fa",
   394 => x"497387e4",
   395 => x"7199ffc3",
   396 => x"fb49c01e",
   397 => x"497387c6",
   398 => x"7129b7c8",
   399 => x"fa49c11e",
   400 => x"86c887fa",
   401 => x"c287c1c6",
   402 => x"4bbff1f7",
   403 => x"87dd029b",
   404 => x"bfdee0c2",
   405 => x"87dec749",
   406 => x"c4059870",
   407 => x"d24bc087",
   408 => x"49e0c287",
   409 => x"c287c3c7",
   410 => x"c658e2e0",
   411 => x"dee0c287",
   412 => x"7378c048",
   413 => x"0599c249",
   414 => x"ebc387ce",
   415 => x"cdd7ff49",
   416 => x"c2497087",
   417 => x"87c20299",
   418 => x"49734cfb",
   419 => x"ce0599c1",
   420 => x"49f4c387",
   421 => x"87f6d6ff",
   422 => x"99c24970",
   423 => x"fa87c202",
   424 => x"c849734c",
   425 => x"87ce0599",
   426 => x"ff49f5c3",
   427 => x"7087dfd6",
   428 => x"0299c249",
   429 => x"f7c287d5",
   430 => x"ca02bff9",
   431 => x"88c14887",
   432 => x"58fdf7c2",
   433 => x"ff87c2c0",
   434 => x"734dc14c",
   435 => x"0599c449",
   436 => x"f2c387ce",
   437 => x"f5d5ff49",
   438 => x"c2497087",
   439 => x"87dc0299",
   440 => x"bff9f7c2",
   441 => x"b7c7487e",
   442 => x"cbc003a8",
   443 => x"c1486e87",
   444 => x"fdf7c280",
   445 => x"87c2c058",
   446 => x"4dc14cfe",
   447 => x"ff49fdc3",
   448 => x"7087cbd5",
   449 => x"0299c249",
   450 => x"c287d5c0",
   451 => x"02bff9f7",
   452 => x"c287c9c0",
   453 => x"c048f9f7",
   454 => x"87c2c078",
   455 => x"4dc14cfd",
   456 => x"ff49fac3",
   457 => x"7087e7d4",
   458 => x"0299c249",
   459 => x"c287d9c0",
   460 => x"48bff9f7",
   461 => x"03a8b7c7",
   462 => x"c287c9c0",
   463 => x"c748f9f7",
   464 => x"87c2c078",
   465 => x"4dc14cfc",
   466 => x"03acb7c0",
   467 => x"c487d1c0",
   468 => x"d8c14a66",
   469 => x"c0026a82",
   470 => x"4b6a87c6",
   471 => x"0f734974",
   472 => x"f0c31ec0",
   473 => x"49dac11e",
   474 => x"c887cef7",
   475 => x"02987086",
   476 => x"c887e2c0",
   477 => x"f7c248a6",
   478 => x"c878bff9",
   479 => x"91cb4966",
   480 => x"714866c4",
   481 => x"6e7e7080",
   482 => x"c8c002bf",
   483 => x"4bbf6e87",
   484 => x"734966c8",
   485 => x"029d750f",
   486 => x"c287c8c0",
   487 => x"49bff9f7",
   488 => x"c287faf2",
   489 => x"02bfe6e0",
   490 => x"4987ddc0",
   491 => x"7087c7c2",
   492 => x"d3c00298",
   493 => x"f9f7c287",
   494 => x"e0f249bf",
   495 => x"f449c087",
   496 => x"e0c287c0",
   497 => x"78c048e6",
   498 => x"daf38ef4",
   499 => x"5b5e0e87",
   500 => x"1e0e5d5c",
   501 => x"f7c24c71",
   502 => x"c149bff5",
   503 => x"c14da1cd",
   504 => x"7e6981d1",
   505 => x"cf029c74",
   506 => x"4ba5c487",
   507 => x"f7c27b74",
   508 => x"f249bff5",
   509 => x"7b6e87f9",
   510 => x"c4059c74",
   511 => x"c24bc087",
   512 => x"734bc187",
   513 => x"87faf249",
   514 => x"c70266d4",
   515 => x"87da4987",
   516 => x"87c24a70",
   517 => x"e0c24ac0",
   518 => x"f2265aea",
   519 => x"000087c9",
   520 => x"00000000",
   521 => x"00000000",
   522 => x"711e0000",
   523 => x"bfc8ff4a",
   524 => x"48a17249",
   525 => x"ff1e4f26",
   526 => x"fe89bfc8",
   527 => x"c0c0c0c0",
   528 => x"c401a9c0",
   529 => x"c24ac087",
   530 => x"724ac187",
   531 => x"1e4f2648",
   532 => x"bfdde2c2",
   533 => x"c2b9c149",
   534 => x"ff59e1e2",
   535 => x"ffc348d4",
   536 => x"48d0ff78",
   537 => x"ff78e1c0",
   538 => x"78c148d4",
   539 => x"787131c4",
   540 => x"c048d0ff",
   541 => x"4f2678e0",
   542 => x"d1e2c21e",
   543 => x"dcf2c21e",
   544 => x"c0fcfd49",
   545 => x"7086c487",
   546 => x"87c30298",
   547 => x"2687c0ff",
   548 => x"4b35314f",
   549 => x"20205a48",
   550 => x"47464320",
   551 => x"00000000",
   552 => x"5b5e0e00",
   553 => x"c20e5d5c",
   554 => x"4abfe9f7",
   555 => x"bfcae4c2",
   556 => x"bc724c49",
   557 => x"c6ff4d71",
   558 => x"4bc087eb",
   559 => x"99d04974",
   560 => x"87e7c002",
   561 => x"c848d0ff",
   562 => x"d4ff78e1",
   563 => x"7578c548",
   564 => x"0299d049",
   565 => x"f0c387c3",
   566 => x"f8e4c278",
   567 => x"11817349",
   568 => x"08d4ff48",
   569 => x"48d0ff78",
   570 => x"c178e0c0",
   571 => x"c8832d2c",
   572 => x"c7ff04ab",
   573 => x"e4c5ff87",
   574 => x"cae4c287",
   575 => x"e9f7c248",
   576 => x"4d2678bf",
   577 => x"4b264c26",
   578 => x"00004f26",
   579 => x"c11e0000",
   580 => x"de48d0e7",
   581 => x"e1e4c250",
   582 => x"f1d9fe49",
   583 => x"2648c087",
   584 => x"4f544a4f",
   585 => x"55525455",
   586 => x"4352414e",
   587 => x"dff21e00",
   588 => x"87edfd87",
   589 => x"4f2687f8",
   590 => x"25261e16",
   591 => x"3e3d362e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
