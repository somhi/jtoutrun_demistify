
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c0",x"f8",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c0",x"f8",x"c2"),
    14 => (x"48",x"c0",x"e5",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ed",x"e5"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"81",x"48",x"73",x"1e"),
    47 => (x"72",x"05",x"a9",x"73"),
    48 => (x"26",x"87",x"f9",x"53"),
    49 => (x"4a",x"71",x"1e",x"4f"),
    50 => (x"48",x"49",x"66",x"c4"),
    51 => (x"a6",x"c8",x"88",x"c1"),
    52 => (x"02",x"99",x"71",x"58"),
    53 => (x"d4",x"ff",x"87",x"d6"),
    54 => (x"78",x"ff",x"c3",x"48"),
    55 => (x"66",x"c4",x"52",x"68"),
    56 => (x"88",x"c1",x"48",x"49"),
    57 => (x"71",x"58",x"a6",x"c8"),
    58 => (x"87",x"ea",x"05",x"99"),
    59 => (x"73",x"1e",x"4f",x"26"),
    60 => (x"4b",x"d4",x"ff",x"1e"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"7b",x"ff",x"c3",x"4a"),
    63 => (x"32",x"c8",x"49",x"6b"),
    64 => (x"ff",x"c3",x"b1",x"72"),
    65 => (x"c8",x"4a",x"6b",x"7b"),
    66 => (x"c3",x"b2",x"71",x"31"),
    67 => (x"49",x"6b",x"7b",x"ff"),
    68 => (x"b1",x"72",x"32",x"c8"),
    69 => (x"87",x"c4",x"48",x"71"),
    70 => (x"4c",x"26",x"4d",x"26"),
    71 => (x"4f",x"26",x"4b",x"26"),
    72 => (x"5c",x"5b",x"5e",x"0e"),
    73 => (x"4a",x"71",x"0e",x"5d"),
    74 => (x"72",x"4c",x"d4",x"ff"),
    75 => (x"99",x"ff",x"c3",x"49"),
    76 => (x"e5",x"c2",x"7c",x"71"),
    77 => (x"c8",x"05",x"bf",x"c0"),
    78 => (x"48",x"66",x"d0",x"87"),
    79 => (x"a6",x"d4",x"30",x"c9"),
    80 => (x"49",x"66",x"d0",x"58"),
    81 => (x"ff",x"c3",x"29",x"d8"),
    82 => (x"d0",x"7c",x"71",x"99"),
    83 => (x"29",x"d0",x"49",x"66"),
    84 => (x"71",x"99",x"ff",x"c3"),
    85 => (x"49",x"66",x"d0",x"7c"),
    86 => (x"ff",x"c3",x"29",x"c8"),
    87 => (x"d0",x"7c",x"71",x"99"),
    88 => (x"ff",x"c3",x"49",x"66"),
    89 => (x"72",x"7c",x"71",x"99"),
    90 => (x"c3",x"29",x"d0",x"49"),
    91 => (x"7c",x"71",x"99",x"ff"),
    92 => (x"f0",x"c9",x"4b",x"6c"),
    93 => (x"ff",x"c3",x"4d",x"ff"),
    94 => (x"87",x"d0",x"05",x"ab"),
    95 => (x"6c",x"7c",x"ff",x"c3"),
    96 => (x"02",x"8d",x"c1",x"4b"),
    97 => (x"ff",x"c3",x"87",x"c6"),
    98 => (x"87",x"f0",x"02",x"ab"),
    99 => (x"c7",x"fe",x"48",x"73"),
   100 => (x"49",x"c0",x"1e",x"87"),
   101 => (x"c3",x"48",x"d4",x"ff"),
   102 => (x"81",x"c1",x"78",x"ff"),
   103 => (x"a9",x"b7",x"c8",x"c3"),
   104 => (x"26",x"87",x"f1",x"04"),
   105 => (x"1e",x"73",x"1e",x"4f"),
   106 => (x"f8",x"c4",x"87",x"e7"),
   107 => (x"1e",x"c0",x"4b",x"df"),
   108 => (x"c1",x"f0",x"ff",x"c0"),
   109 => (x"e7",x"fd",x"49",x"f7"),
   110 => (x"c1",x"86",x"c4",x"87"),
   111 => (x"ea",x"c0",x"05",x"a8"),
   112 => (x"48",x"d4",x"ff",x"87"),
   113 => (x"c1",x"78",x"ff",x"c3"),
   114 => (x"c0",x"c0",x"c0",x"c0"),
   115 => (x"e1",x"c0",x"1e",x"c0"),
   116 => (x"49",x"e9",x"c1",x"f0"),
   117 => (x"c4",x"87",x"c9",x"fd"),
   118 => (x"05",x"98",x"70",x"86"),
   119 => (x"d4",x"ff",x"87",x"ca"),
   120 => (x"78",x"ff",x"c3",x"48"),
   121 => (x"87",x"cb",x"48",x"c1"),
   122 => (x"c1",x"87",x"e6",x"fe"),
   123 => (x"fd",x"fe",x"05",x"8b"),
   124 => (x"fc",x"48",x"c0",x"87"),
   125 => (x"73",x"1e",x"87",x"e6"),
   126 => (x"48",x"d4",x"ff",x"1e"),
   127 => (x"d3",x"78",x"ff",x"c3"),
   128 => (x"c0",x"1e",x"c0",x"4b"),
   129 => (x"c1",x"c1",x"f0",x"ff"),
   130 => (x"87",x"d4",x"fc",x"49"),
   131 => (x"98",x"70",x"86",x"c4"),
   132 => (x"ff",x"87",x"ca",x"05"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"cb",x"48",x"c1",x"78"),
   135 => (x"87",x"f1",x"fd",x"87"),
   136 => (x"ff",x"05",x"8b",x"c1"),
   137 => (x"48",x"c0",x"87",x"db"),
   138 => (x"0e",x"87",x"f1",x"fb"),
   139 => (x"0e",x"5c",x"5b",x"5e"),
   140 => (x"fd",x"4c",x"d4",x"ff"),
   141 => (x"ea",x"c6",x"87",x"db"),
   142 => (x"f0",x"e1",x"c0",x"1e"),
   143 => (x"fb",x"49",x"c8",x"c1"),
   144 => (x"86",x"c4",x"87",x"de"),
   145 => (x"c8",x"02",x"a8",x"c1"),
   146 => (x"87",x"ea",x"fe",x"87"),
   147 => (x"e2",x"c1",x"48",x"c0"),
   148 => (x"87",x"da",x"fa",x"87"),
   149 => (x"ff",x"cf",x"49",x"70"),
   150 => (x"ea",x"c6",x"99",x"ff"),
   151 => (x"87",x"c8",x"02",x"a9"),
   152 => (x"c0",x"87",x"d3",x"fe"),
   153 => (x"87",x"cb",x"c1",x"48"),
   154 => (x"c0",x"7c",x"ff",x"c3"),
   155 => (x"f4",x"fc",x"4b",x"f1"),
   156 => (x"02",x"98",x"70",x"87"),
   157 => (x"c0",x"87",x"eb",x"c0"),
   158 => (x"f0",x"ff",x"c0",x"1e"),
   159 => (x"fa",x"49",x"fa",x"c1"),
   160 => (x"86",x"c4",x"87",x"de"),
   161 => (x"d9",x"05",x"98",x"70"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"ff",x"c3",x"49",x"6c"),
   164 => (x"7c",x"7c",x"7c",x"7c"),
   165 => (x"02",x"99",x"c0",x"c1"),
   166 => (x"48",x"c1",x"87",x"c4"),
   167 => (x"48",x"c0",x"87",x"d5"),
   168 => (x"ab",x"c2",x"87",x"d1"),
   169 => (x"c0",x"87",x"c4",x"05"),
   170 => (x"c1",x"87",x"c8",x"48"),
   171 => (x"fd",x"fe",x"05",x"8b"),
   172 => (x"f9",x"48",x"c0",x"87"),
   173 => (x"73",x"1e",x"87",x"e4"),
   174 => (x"c0",x"e5",x"c2",x"1e"),
   175 => (x"c7",x"78",x"c1",x"48"),
   176 => (x"48",x"d0",x"ff",x"4b"),
   177 => (x"c8",x"fb",x"78",x"c2"),
   178 => (x"48",x"d0",x"ff",x"87"),
   179 => (x"1e",x"c0",x"78",x"c3"),
   180 => (x"c1",x"d0",x"e5",x"c0"),
   181 => (x"c7",x"f9",x"49",x"c0"),
   182 => (x"c1",x"86",x"c4",x"87"),
   183 => (x"87",x"c1",x"05",x"a8"),
   184 => (x"05",x"ab",x"c2",x"4b"),
   185 => (x"48",x"c0",x"87",x"c5"),
   186 => (x"c1",x"87",x"f9",x"c0"),
   187 => (x"d0",x"ff",x"05",x"8b"),
   188 => (x"87",x"f7",x"fc",x"87"),
   189 => (x"58",x"c4",x"e5",x"c2"),
   190 => (x"cd",x"05",x"98",x"70"),
   191 => (x"c0",x"1e",x"c1",x"87"),
   192 => (x"d0",x"c1",x"f0",x"ff"),
   193 => (x"87",x"d8",x"f8",x"49"),
   194 => (x"d4",x"ff",x"86",x"c4"),
   195 => (x"78",x"ff",x"c3",x"48"),
   196 => (x"c2",x"87",x"fc",x"c2"),
   197 => (x"ff",x"58",x"c8",x"e5"),
   198 => (x"78",x"c2",x"48",x"d0"),
   199 => (x"c3",x"48",x"d4",x"ff"),
   200 => (x"48",x"c1",x"78",x"ff"),
   201 => (x"0e",x"87",x"f5",x"f7"),
   202 => (x"5d",x"5c",x"5b",x"5e"),
   203 => (x"c0",x"4b",x"71",x"0e"),
   204 => (x"cd",x"ee",x"c5",x"4c"),
   205 => (x"d4",x"ff",x"4a",x"df"),
   206 => (x"78",x"ff",x"c3",x"48"),
   207 => (x"fe",x"c3",x"49",x"68"),
   208 => (x"fd",x"c0",x"05",x"a9"),
   209 => (x"73",x"4d",x"70",x"87"),
   210 => (x"87",x"cc",x"02",x"9b"),
   211 => (x"73",x"1e",x"66",x"d0"),
   212 => (x"87",x"f1",x"f5",x"49"),
   213 => (x"87",x"d6",x"86",x"c4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"ff",x"c3",x"78",x"d1"),
   216 => (x"48",x"66",x"d0",x"7d"),
   217 => (x"a6",x"d4",x"88",x"c1"),
   218 => (x"05",x"98",x"70",x"58"),
   219 => (x"d4",x"ff",x"87",x"f0"),
   220 => (x"78",x"ff",x"c3",x"48"),
   221 => (x"05",x"9b",x"73",x"78"),
   222 => (x"d0",x"ff",x"87",x"c5"),
   223 => (x"c1",x"78",x"d0",x"48"),
   224 => (x"8a",x"c1",x"4c",x"4a"),
   225 => (x"87",x"ee",x"fe",x"05"),
   226 => (x"cb",x"f6",x"48",x"74"),
   227 => (x"1e",x"73",x"1e",x"87"),
   228 => (x"4b",x"c0",x"4a",x"71"),
   229 => (x"c3",x"48",x"d4",x"ff"),
   230 => (x"d0",x"ff",x"78",x"ff"),
   231 => (x"78",x"c3",x"c4",x"48"),
   232 => (x"c3",x"48",x"d4",x"ff"),
   233 => (x"1e",x"72",x"78",x"ff"),
   234 => (x"c1",x"f0",x"ff",x"c0"),
   235 => (x"ef",x"f5",x"49",x"d1"),
   236 => (x"70",x"86",x"c4",x"87"),
   237 => (x"87",x"d2",x"05",x"98"),
   238 => (x"cc",x"1e",x"c0",x"c8"),
   239 => (x"e6",x"fd",x"49",x"66"),
   240 => (x"70",x"86",x"c4",x"87"),
   241 => (x"48",x"d0",x"ff",x"4b"),
   242 => (x"48",x"73",x"78",x"c2"),
   243 => (x"0e",x"87",x"cd",x"f5"),
   244 => (x"5d",x"5c",x"5b",x"5e"),
   245 => (x"c0",x"1e",x"c0",x"0e"),
   246 => (x"c9",x"c1",x"f0",x"ff"),
   247 => (x"87",x"c0",x"f5",x"49"),
   248 => (x"e5",x"c2",x"1e",x"d2"),
   249 => (x"fe",x"fc",x"49",x"c8"),
   250 => (x"c0",x"86",x"c8",x"87"),
   251 => (x"d2",x"84",x"c1",x"4c"),
   252 => (x"f8",x"04",x"ac",x"b7"),
   253 => (x"c8",x"e5",x"c2",x"87"),
   254 => (x"c3",x"49",x"bf",x"97"),
   255 => (x"c0",x"c1",x"99",x"c0"),
   256 => (x"e7",x"c0",x"05",x"a9"),
   257 => (x"cf",x"e5",x"c2",x"87"),
   258 => (x"d0",x"49",x"bf",x"97"),
   259 => (x"d0",x"e5",x"c2",x"31"),
   260 => (x"c8",x"4a",x"bf",x"97"),
   261 => (x"c2",x"b1",x"72",x"32"),
   262 => (x"bf",x"97",x"d1",x"e5"),
   263 => (x"4c",x"71",x"b1",x"4a"),
   264 => (x"ff",x"ff",x"ff",x"cf"),
   265 => (x"ca",x"84",x"c1",x"9c"),
   266 => (x"87",x"e7",x"c1",x"34"),
   267 => (x"97",x"d1",x"e5",x"c2"),
   268 => (x"31",x"c1",x"49",x"bf"),
   269 => (x"e5",x"c2",x"99",x"c6"),
   270 => (x"4a",x"bf",x"97",x"d2"),
   271 => (x"72",x"2a",x"b7",x"c7"),
   272 => (x"cd",x"e5",x"c2",x"b1"),
   273 => (x"4d",x"4a",x"bf",x"97"),
   274 => (x"e5",x"c2",x"9d",x"cf"),
   275 => (x"4a",x"bf",x"97",x"ce"),
   276 => (x"32",x"ca",x"9a",x"c3"),
   277 => (x"97",x"cf",x"e5",x"c2"),
   278 => (x"33",x"c2",x"4b",x"bf"),
   279 => (x"e5",x"c2",x"b2",x"73"),
   280 => (x"4b",x"bf",x"97",x"d0"),
   281 => (x"c6",x"9b",x"c0",x"c3"),
   282 => (x"b2",x"73",x"2b",x"b7"),
   283 => (x"48",x"c1",x"81",x"c2"),
   284 => (x"49",x"70",x"30",x"71"),
   285 => (x"30",x"75",x"48",x"c1"),
   286 => (x"4c",x"72",x"4d",x"70"),
   287 => (x"94",x"71",x"84",x"c1"),
   288 => (x"ad",x"b7",x"c0",x"c8"),
   289 => (x"c1",x"87",x"cc",x"06"),
   290 => (x"c8",x"2d",x"b7",x"34"),
   291 => (x"01",x"ad",x"b7",x"c0"),
   292 => (x"74",x"87",x"f4",x"ff"),
   293 => (x"87",x"c0",x"f2",x"48"),
   294 => (x"5c",x"5b",x"5e",x"0e"),
   295 => (x"86",x"f8",x"0e",x"5d"),
   296 => (x"48",x"ee",x"ed",x"c2"),
   297 => (x"e5",x"c2",x"78",x"c0"),
   298 => (x"49",x"c0",x"1e",x"e6"),
   299 => (x"c4",x"87",x"de",x"fb"),
   300 => (x"05",x"98",x"70",x"86"),
   301 => (x"48",x"c0",x"87",x"c5"),
   302 => (x"c0",x"87",x"ce",x"c9"),
   303 => (x"c0",x"7e",x"c1",x"4d"),
   304 => (x"49",x"bf",x"d8",x"f5"),
   305 => (x"4a",x"dc",x"e6",x"c2"),
   306 => (x"ee",x"4b",x"c8",x"71"),
   307 => (x"98",x"70",x"87",x"dc"),
   308 => (x"c0",x"87",x"c2",x"05"),
   309 => (x"d4",x"f5",x"c0",x"7e"),
   310 => (x"e6",x"c2",x"49",x"bf"),
   311 => (x"c8",x"71",x"4a",x"f8"),
   312 => (x"87",x"c6",x"ee",x"4b"),
   313 => (x"c2",x"05",x"98",x"70"),
   314 => (x"6e",x"7e",x"c0",x"87"),
   315 => (x"87",x"fd",x"c0",x"02"),
   316 => (x"bf",x"ec",x"ec",x"c2"),
   317 => (x"e4",x"ed",x"c2",x"4d"),
   318 => (x"48",x"7e",x"bf",x"9f"),
   319 => (x"a8",x"ea",x"d6",x"c5"),
   320 => (x"c2",x"87",x"c7",x"05"),
   321 => (x"4d",x"bf",x"ec",x"ec"),
   322 => (x"48",x"6e",x"87",x"ce"),
   323 => (x"a8",x"d5",x"e9",x"ca"),
   324 => (x"c0",x"87",x"c5",x"02"),
   325 => (x"87",x"f1",x"c7",x"48"),
   326 => (x"1e",x"e6",x"e5",x"c2"),
   327 => (x"ec",x"f9",x"49",x"75"),
   328 => (x"70",x"86",x"c4",x"87"),
   329 => (x"87",x"c5",x"05",x"98"),
   330 => (x"dc",x"c7",x"48",x"c0"),
   331 => (x"d4",x"f5",x"c0",x"87"),
   332 => (x"e6",x"c2",x"49",x"bf"),
   333 => (x"c8",x"71",x"4a",x"f8"),
   334 => (x"87",x"ee",x"ec",x"4b"),
   335 => (x"c8",x"05",x"98",x"70"),
   336 => (x"ee",x"ed",x"c2",x"87"),
   337 => (x"da",x"78",x"c1",x"48"),
   338 => (x"d8",x"f5",x"c0",x"87"),
   339 => (x"e6",x"c2",x"49",x"bf"),
   340 => (x"c8",x"71",x"4a",x"dc"),
   341 => (x"87",x"d2",x"ec",x"4b"),
   342 => (x"c0",x"02",x"98",x"70"),
   343 => (x"48",x"c0",x"87",x"c5"),
   344 => (x"c2",x"87",x"e6",x"c6"),
   345 => (x"bf",x"97",x"e4",x"ed"),
   346 => (x"a9",x"d5",x"c1",x"49"),
   347 => (x"87",x"cd",x"c0",x"05"),
   348 => (x"97",x"e5",x"ed",x"c2"),
   349 => (x"ea",x"c2",x"49",x"bf"),
   350 => (x"c5",x"c0",x"02",x"a9"),
   351 => (x"c6",x"48",x"c0",x"87"),
   352 => (x"e5",x"c2",x"87",x"c7"),
   353 => (x"7e",x"bf",x"97",x"e6"),
   354 => (x"a8",x"e9",x"c3",x"48"),
   355 => (x"87",x"ce",x"c0",x"02"),
   356 => (x"eb",x"c3",x"48",x"6e"),
   357 => (x"c5",x"c0",x"02",x"a8"),
   358 => (x"c5",x"48",x"c0",x"87"),
   359 => (x"e5",x"c2",x"87",x"eb"),
   360 => (x"49",x"bf",x"97",x"f1"),
   361 => (x"cc",x"c0",x"05",x"99"),
   362 => (x"f2",x"e5",x"c2",x"87"),
   363 => (x"c2",x"49",x"bf",x"97"),
   364 => (x"c5",x"c0",x"02",x"a9"),
   365 => (x"c5",x"48",x"c0",x"87"),
   366 => (x"e5",x"c2",x"87",x"cf"),
   367 => (x"48",x"bf",x"97",x"f3"),
   368 => (x"58",x"ea",x"ed",x"c2"),
   369 => (x"c1",x"48",x"4c",x"70"),
   370 => (x"ee",x"ed",x"c2",x"88"),
   371 => (x"f4",x"e5",x"c2",x"58"),
   372 => (x"75",x"49",x"bf",x"97"),
   373 => (x"f5",x"e5",x"c2",x"81"),
   374 => (x"c8",x"4a",x"bf",x"97"),
   375 => (x"7e",x"a1",x"72",x"32"),
   376 => (x"48",x"fb",x"f1",x"c2"),
   377 => (x"e5",x"c2",x"78",x"6e"),
   378 => (x"48",x"bf",x"97",x"f6"),
   379 => (x"c2",x"58",x"a6",x"c8"),
   380 => (x"02",x"bf",x"ee",x"ed"),
   381 => (x"c0",x"87",x"d4",x"c2"),
   382 => (x"49",x"bf",x"d4",x"f5"),
   383 => (x"4a",x"f8",x"e6",x"c2"),
   384 => (x"e9",x"4b",x"c8",x"71"),
   385 => (x"98",x"70",x"87",x"e4"),
   386 => (x"87",x"c5",x"c0",x"02"),
   387 => (x"f8",x"c3",x"48",x"c0"),
   388 => (x"e6",x"ed",x"c2",x"87"),
   389 => (x"f2",x"c2",x"4c",x"bf"),
   390 => (x"e6",x"c2",x"5c",x"cf"),
   391 => (x"49",x"bf",x"97",x"cb"),
   392 => (x"e6",x"c2",x"31",x"c8"),
   393 => (x"4a",x"bf",x"97",x"ca"),
   394 => (x"e6",x"c2",x"49",x"a1"),
   395 => (x"4a",x"bf",x"97",x"cc"),
   396 => (x"a1",x"72",x"32",x"d0"),
   397 => (x"cd",x"e6",x"c2",x"49"),
   398 => (x"d8",x"4a",x"bf",x"97"),
   399 => (x"49",x"a1",x"72",x"32"),
   400 => (x"c2",x"91",x"66",x"c4"),
   401 => (x"81",x"bf",x"fb",x"f1"),
   402 => (x"59",x"c3",x"f2",x"c2"),
   403 => (x"97",x"d3",x"e6",x"c2"),
   404 => (x"32",x"c8",x"4a",x"bf"),
   405 => (x"97",x"d2",x"e6",x"c2"),
   406 => (x"4a",x"a2",x"4b",x"bf"),
   407 => (x"97",x"d4",x"e6",x"c2"),
   408 => (x"33",x"d0",x"4b",x"bf"),
   409 => (x"c2",x"4a",x"a2",x"73"),
   410 => (x"bf",x"97",x"d5",x"e6"),
   411 => (x"d8",x"9b",x"cf",x"4b"),
   412 => (x"4a",x"a2",x"73",x"33"),
   413 => (x"5a",x"c7",x"f2",x"c2"),
   414 => (x"bf",x"c3",x"f2",x"c2"),
   415 => (x"74",x"8a",x"c2",x"4a"),
   416 => (x"c7",x"f2",x"c2",x"92"),
   417 => (x"78",x"a1",x"72",x"48"),
   418 => (x"c2",x"87",x"ca",x"c1"),
   419 => (x"bf",x"97",x"f8",x"e5"),
   420 => (x"c2",x"31",x"c8",x"49"),
   421 => (x"bf",x"97",x"f7",x"e5"),
   422 => (x"c2",x"49",x"a1",x"4a"),
   423 => (x"c2",x"59",x"f6",x"ed"),
   424 => (x"49",x"bf",x"f2",x"ed"),
   425 => (x"ff",x"c7",x"31",x"c5"),
   426 => (x"c2",x"29",x"c9",x"81"),
   427 => (x"c2",x"59",x"cf",x"f2"),
   428 => (x"bf",x"97",x"fd",x"e5"),
   429 => (x"c2",x"32",x"c8",x"4a"),
   430 => (x"bf",x"97",x"fc",x"e5"),
   431 => (x"c4",x"4a",x"a2",x"4b"),
   432 => (x"82",x"6e",x"92",x"66"),
   433 => (x"5a",x"cb",x"f2",x"c2"),
   434 => (x"48",x"c3",x"f2",x"c2"),
   435 => (x"f1",x"c2",x"78",x"c0"),
   436 => (x"a1",x"72",x"48",x"ff"),
   437 => (x"cf",x"f2",x"c2",x"78"),
   438 => (x"c3",x"f2",x"c2",x"48"),
   439 => (x"f2",x"c2",x"78",x"bf"),
   440 => (x"f2",x"c2",x"48",x"d3"),
   441 => (x"c2",x"78",x"bf",x"c7"),
   442 => (x"02",x"bf",x"ee",x"ed"),
   443 => (x"74",x"87",x"c9",x"c0"),
   444 => (x"70",x"30",x"c4",x"48"),
   445 => (x"87",x"c9",x"c0",x"7e"),
   446 => (x"bf",x"cb",x"f2",x"c2"),
   447 => (x"70",x"30",x"c4",x"48"),
   448 => (x"f2",x"ed",x"c2",x"7e"),
   449 => (x"c1",x"78",x"6e",x"48"),
   450 => (x"26",x"8e",x"f8",x"48"),
   451 => (x"26",x"4c",x"26",x"4d"),
   452 => (x"0e",x"4f",x"26",x"4b"),
   453 => (x"5d",x"5c",x"5b",x"5e"),
   454 => (x"c2",x"4a",x"71",x"0e"),
   455 => (x"02",x"bf",x"ee",x"ed"),
   456 => (x"4b",x"72",x"87",x"cb"),
   457 => (x"4c",x"72",x"2b",x"c7"),
   458 => (x"c9",x"9c",x"ff",x"c1"),
   459 => (x"c8",x"4b",x"72",x"87"),
   460 => (x"c3",x"4c",x"72",x"2b"),
   461 => (x"f1",x"c2",x"9c",x"ff"),
   462 => (x"c0",x"83",x"bf",x"fb"),
   463 => (x"ab",x"bf",x"d0",x"f5"),
   464 => (x"c0",x"87",x"d9",x"02"),
   465 => (x"c2",x"5b",x"d4",x"f5"),
   466 => (x"73",x"1e",x"e6",x"e5"),
   467 => (x"87",x"fd",x"f0",x"49"),
   468 => (x"98",x"70",x"86",x"c4"),
   469 => (x"c0",x"87",x"c5",x"05"),
   470 => (x"87",x"e6",x"c0",x"48"),
   471 => (x"bf",x"ee",x"ed",x"c2"),
   472 => (x"74",x"87",x"d2",x"02"),
   473 => (x"c2",x"91",x"c4",x"49"),
   474 => (x"69",x"81",x"e6",x"e5"),
   475 => (x"ff",x"ff",x"cf",x"4d"),
   476 => (x"cb",x"9d",x"ff",x"ff"),
   477 => (x"c2",x"49",x"74",x"87"),
   478 => (x"e6",x"e5",x"c2",x"91"),
   479 => (x"4d",x"69",x"9f",x"81"),
   480 => (x"c6",x"fe",x"48",x"75"),
   481 => (x"5b",x"5e",x"0e",x"87"),
   482 => (x"f8",x"0e",x"5d",x"5c"),
   483 => (x"9c",x"4c",x"71",x"86"),
   484 => (x"c0",x"87",x"c5",x"05"),
   485 => (x"87",x"c1",x"c3",x"48"),
   486 => (x"6e",x"7e",x"a4",x"c8"),
   487 => (x"d8",x"78",x"c0",x"48"),
   488 => (x"87",x"c7",x"02",x"66"),
   489 => (x"bf",x"97",x"66",x"d8"),
   490 => (x"c0",x"87",x"c5",x"05"),
   491 => (x"87",x"e9",x"c2",x"48"),
   492 => (x"49",x"c1",x"1e",x"c0"),
   493 => (x"c4",x"87",x"fd",x"ce"),
   494 => (x"9d",x"4d",x"70",x"86"),
   495 => (x"87",x"c2",x"c1",x"02"),
   496 => (x"4a",x"f6",x"ed",x"c2"),
   497 => (x"e2",x"49",x"66",x"d8"),
   498 => (x"98",x"70",x"87",x"c5"),
   499 => (x"87",x"f2",x"c0",x"02"),
   500 => (x"66",x"d8",x"4a",x"75"),
   501 => (x"e2",x"4b",x"cb",x"49"),
   502 => (x"98",x"70",x"87",x"ea"),
   503 => (x"87",x"e2",x"c0",x"02"),
   504 => (x"9d",x"75",x"1e",x"c0"),
   505 => (x"c8",x"87",x"c7",x"02"),
   506 => (x"78",x"c0",x"48",x"a6"),
   507 => (x"a6",x"c8",x"87",x"c5"),
   508 => (x"c8",x"78",x"c1",x"48"),
   509 => (x"fb",x"cd",x"49",x"66"),
   510 => (x"70",x"86",x"c4",x"87"),
   511 => (x"fe",x"05",x"9d",x"4d"),
   512 => (x"9d",x"75",x"87",x"fe"),
   513 => (x"87",x"cf",x"c1",x"02"),
   514 => (x"6e",x"49",x"a5",x"dc"),
   515 => (x"da",x"78",x"69",x"48"),
   516 => (x"a6",x"c4",x"49",x"a5"),
   517 => (x"78",x"a4",x"c4",x"48"),
   518 => (x"c4",x"48",x"69",x"9f"),
   519 => (x"c2",x"78",x"08",x"66"),
   520 => (x"02",x"bf",x"ee",x"ed"),
   521 => (x"a5",x"d4",x"87",x"d2"),
   522 => (x"49",x"69",x"9f",x"49"),
   523 => (x"99",x"ff",x"ff",x"c0"),
   524 => (x"30",x"d0",x"48",x"71"),
   525 => (x"87",x"c2",x"7e",x"70"),
   526 => (x"49",x"6e",x"7e",x"c0"),
   527 => (x"bf",x"66",x"c4",x"48"),
   528 => (x"08",x"66",x"c4",x"80"),
   529 => (x"cc",x"7c",x"c0",x"78"),
   530 => (x"66",x"c4",x"49",x"a4"),
   531 => (x"a4",x"d0",x"79",x"bf"),
   532 => (x"c1",x"79",x"c0",x"49"),
   533 => (x"c0",x"87",x"c2",x"48"),
   534 => (x"fa",x"8e",x"f8",x"48"),
   535 => (x"5e",x"0e",x"87",x"ed"),
   536 => (x"0e",x"5d",x"5c",x"5b"),
   537 => (x"02",x"9c",x"4c",x"71"),
   538 => (x"c8",x"87",x"ca",x"c1"),
   539 => (x"02",x"69",x"49",x"a4"),
   540 => (x"d0",x"87",x"c2",x"c1"),
   541 => (x"49",x"6c",x"4a",x"66"),
   542 => (x"5a",x"a6",x"d4",x"82"),
   543 => (x"b9",x"4d",x"66",x"d0"),
   544 => (x"bf",x"ea",x"ed",x"c2"),
   545 => (x"72",x"ba",x"ff",x"4a"),
   546 => (x"02",x"99",x"71",x"99"),
   547 => (x"c4",x"87",x"e4",x"c0"),
   548 => (x"49",x"6b",x"4b",x"a4"),
   549 => (x"70",x"87",x"fc",x"f9"),
   550 => (x"e6",x"ed",x"c2",x"7b"),
   551 => (x"81",x"6c",x"49",x"bf"),
   552 => (x"b9",x"75",x"7c",x"71"),
   553 => (x"bf",x"ea",x"ed",x"c2"),
   554 => (x"72",x"ba",x"ff",x"4a"),
   555 => (x"05",x"99",x"71",x"99"),
   556 => (x"75",x"87",x"dc",x"ff"),
   557 => (x"87",x"d3",x"f9",x"7c"),
   558 => (x"71",x"1e",x"73",x"1e"),
   559 => (x"c7",x"02",x"9b",x"4b"),
   560 => (x"49",x"a3",x"c8",x"87"),
   561 => (x"87",x"c5",x"05",x"69"),
   562 => (x"f7",x"c0",x"48",x"c0"),
   563 => (x"ff",x"f1",x"c2",x"87"),
   564 => (x"a3",x"c4",x"4a",x"bf"),
   565 => (x"c2",x"49",x"69",x"49"),
   566 => (x"e6",x"ed",x"c2",x"89"),
   567 => (x"a2",x"71",x"91",x"bf"),
   568 => (x"ea",x"ed",x"c2",x"4a"),
   569 => (x"99",x"6b",x"49",x"bf"),
   570 => (x"c0",x"4a",x"a2",x"71"),
   571 => (x"c8",x"5a",x"d4",x"f5"),
   572 => (x"49",x"72",x"1e",x"66"),
   573 => (x"c4",x"87",x"d6",x"ea"),
   574 => (x"05",x"98",x"70",x"86"),
   575 => (x"48",x"c0",x"87",x"c4"),
   576 => (x"48",x"c1",x"87",x"c2"),
   577 => (x"0e",x"87",x"c8",x"f8"),
   578 => (x"0e",x"5c",x"5b",x"5e"),
   579 => (x"d0",x"4b",x"71",x"1e"),
   580 => (x"2c",x"c9",x"4c",x"66"),
   581 => (x"c1",x"02",x"9b",x"73"),
   582 => (x"a3",x"c8",x"87",x"d4"),
   583 => (x"c1",x"02",x"69",x"49"),
   584 => (x"ed",x"c2",x"87",x"cc"),
   585 => (x"ff",x"49",x"bf",x"ea"),
   586 => (x"99",x"4a",x"6b",x"b9"),
   587 => (x"03",x"ac",x"71",x"7e"),
   588 => (x"7b",x"c0",x"87",x"d1"),
   589 => (x"c0",x"49",x"a3",x"d0"),
   590 => (x"4a",x"a3",x"cc",x"79"),
   591 => (x"6a",x"49",x"a3",x"c4"),
   592 => (x"72",x"87",x"c2",x"79"),
   593 => (x"02",x"9c",x"74",x"8c"),
   594 => (x"49",x"87",x"e3",x"c0"),
   595 => (x"fc",x"49",x"73",x"1e"),
   596 => (x"86",x"c4",x"87",x"cc"),
   597 => (x"c7",x"49",x"66",x"d0"),
   598 => (x"cb",x"02",x"99",x"ff"),
   599 => (x"e6",x"e5",x"c2",x"87"),
   600 => (x"fd",x"49",x"73",x"1e"),
   601 => (x"86",x"c4",x"87",x"d2"),
   602 => (x"d0",x"49",x"a3",x"d0"),
   603 => (x"f6",x"26",x"79",x"66"),
   604 => (x"5e",x"0e",x"87",x"db"),
   605 => (x"0e",x"5d",x"5c",x"5b"),
   606 => (x"a6",x"d0",x"86",x"f0"),
   607 => (x"66",x"e4",x"c0",x"59"),
   608 => (x"02",x"66",x"cc",x"4b"),
   609 => (x"c8",x"48",x"87",x"ca"),
   610 => (x"6e",x"7e",x"70",x"80"),
   611 => (x"87",x"c5",x"05",x"bf"),
   612 => (x"ec",x"c3",x"48",x"c0"),
   613 => (x"4c",x"66",x"cc",x"87"),
   614 => (x"49",x"73",x"84",x"d0"),
   615 => (x"6c",x"48",x"a6",x"c4"),
   616 => (x"81",x"66",x"c4",x"78"),
   617 => (x"bf",x"6e",x"80",x"c4"),
   618 => (x"a9",x"66",x"c8",x"78"),
   619 => (x"49",x"87",x"c6",x"06"),
   620 => (x"71",x"89",x"66",x"c4"),
   621 => (x"ab",x"b7",x"c0",x"4b"),
   622 => (x"48",x"87",x"c4",x"01"),
   623 => (x"c4",x"87",x"c2",x"c3"),
   624 => (x"ff",x"c7",x"48",x"66"),
   625 => (x"6e",x"7e",x"70",x"98"),
   626 => (x"87",x"c9",x"c1",x"02"),
   627 => (x"6e",x"49",x"c0",x"c8"),
   628 => (x"c2",x"4a",x"71",x"89"),
   629 => (x"6e",x"4d",x"e6",x"e5"),
   630 => (x"aa",x"b7",x"73",x"85"),
   631 => (x"4a",x"87",x"c1",x"06"),
   632 => (x"c4",x"48",x"49",x"72"),
   633 => (x"7c",x"70",x"80",x"66"),
   634 => (x"c1",x"49",x"8b",x"72"),
   635 => (x"02",x"99",x"71",x"8a"),
   636 => (x"e0",x"c0",x"87",x"d9"),
   637 => (x"50",x"15",x"48",x"66"),
   638 => (x"48",x"66",x"e0",x"c0"),
   639 => (x"e4",x"c0",x"80",x"c1"),
   640 => (x"49",x"72",x"58",x"a6"),
   641 => (x"99",x"71",x"8a",x"c1"),
   642 => (x"c1",x"87",x"e7",x"05"),
   643 => (x"49",x"66",x"d0",x"1e"),
   644 => (x"c4",x"87",x"cb",x"f9"),
   645 => (x"ab",x"b7",x"c0",x"86"),
   646 => (x"87",x"e3",x"c1",x"06"),
   647 => (x"4d",x"66",x"e0",x"c0"),
   648 => (x"ab",x"b7",x"ff",x"c7"),
   649 => (x"87",x"e2",x"c0",x"06"),
   650 => (x"66",x"d0",x"1e",x"75"),
   651 => (x"87",x"c8",x"fa",x"49"),
   652 => (x"6c",x"85",x"c0",x"c8"),
   653 => (x"80",x"c0",x"c8",x"48"),
   654 => (x"c0",x"c8",x"7c",x"70"),
   655 => (x"d4",x"1e",x"c1",x"8b"),
   656 => (x"d9",x"f8",x"49",x"66"),
   657 => (x"c0",x"86",x"c8",x"87"),
   658 => (x"e5",x"c2",x"87",x"ee"),
   659 => (x"66",x"d0",x"1e",x"e6"),
   660 => (x"87",x"e4",x"f9",x"49"),
   661 => (x"e5",x"c2",x"86",x"c4"),
   662 => (x"49",x"73",x"4a",x"e6"),
   663 => (x"70",x"80",x"6c",x"48"),
   664 => (x"c1",x"49",x"73",x"7c"),
   665 => (x"02",x"99",x"71",x"8b"),
   666 => (x"97",x"12",x"87",x"ce"),
   667 => (x"73",x"85",x"c1",x"7d"),
   668 => (x"71",x"8b",x"c1",x"49"),
   669 => (x"87",x"f2",x"05",x"99"),
   670 => (x"01",x"ab",x"b7",x"c0"),
   671 => (x"c1",x"87",x"e1",x"fe"),
   672 => (x"f2",x"8e",x"f0",x"48"),
   673 => (x"5e",x"0e",x"87",x"c5"),
   674 => (x"0e",x"5d",x"5c",x"5b"),
   675 => (x"02",x"9b",x"4b",x"71"),
   676 => (x"a3",x"c8",x"87",x"c7"),
   677 => (x"c5",x"05",x"6d",x"4d"),
   678 => (x"c0",x"48",x"ff",x"87"),
   679 => (x"a3",x"d0",x"87",x"fd"),
   680 => (x"c7",x"49",x"6c",x"4c"),
   681 => (x"d8",x"05",x"99",x"ff"),
   682 => (x"c9",x"02",x"6c",x"87"),
   683 => (x"73",x"1e",x"c1",x"87"),
   684 => (x"87",x"ea",x"f6",x"49"),
   685 => (x"e5",x"c2",x"86",x"c4"),
   686 => (x"49",x"73",x"1e",x"e6"),
   687 => (x"c4",x"87",x"f9",x"f7"),
   688 => (x"6d",x"4a",x"6c",x"86"),
   689 => (x"87",x"c4",x"04",x"aa"),
   690 => (x"87",x"cf",x"48",x"ff"),
   691 => (x"72",x"7c",x"a2",x"c1"),
   692 => (x"99",x"ff",x"c7",x"49"),
   693 => (x"81",x"e6",x"e5",x"c2"),
   694 => (x"f0",x"48",x"69",x"97"),
   695 => (x"73",x"1e",x"87",x"ed"),
   696 => (x"9b",x"4b",x"71",x"1e"),
   697 => (x"87",x"e4",x"c0",x"02"),
   698 => (x"5b",x"d3",x"f2",x"c2"),
   699 => (x"8a",x"c2",x"4a",x"73"),
   700 => (x"bf",x"e6",x"ed",x"c2"),
   701 => (x"f1",x"c2",x"92",x"49"),
   702 => (x"72",x"48",x"bf",x"ff"),
   703 => (x"d7",x"f2",x"c2",x"80"),
   704 => (x"c4",x"48",x"71",x"58"),
   705 => (x"f6",x"ed",x"c2",x"30"),
   706 => (x"87",x"ed",x"c0",x"58"),
   707 => (x"48",x"cf",x"f2",x"c2"),
   708 => (x"bf",x"c3",x"f2",x"c2"),
   709 => (x"d3",x"f2",x"c2",x"78"),
   710 => (x"c7",x"f2",x"c2",x"48"),
   711 => (x"ed",x"c2",x"78",x"bf"),
   712 => (x"c9",x"02",x"bf",x"ee"),
   713 => (x"e6",x"ed",x"c2",x"87"),
   714 => (x"31",x"c4",x"49",x"bf"),
   715 => (x"f2",x"c2",x"87",x"c7"),
   716 => (x"c4",x"49",x"bf",x"cb"),
   717 => (x"f6",x"ed",x"c2",x"31"),
   718 => (x"87",x"d3",x"ef",x"59"),
   719 => (x"5c",x"5b",x"5e",x"0e"),
   720 => (x"c0",x"4a",x"71",x"0e"),
   721 => (x"02",x"9a",x"72",x"4b"),
   722 => (x"da",x"87",x"e1",x"c0"),
   723 => (x"69",x"9f",x"49",x"a2"),
   724 => (x"ee",x"ed",x"c2",x"4b"),
   725 => (x"87",x"cf",x"02",x"bf"),
   726 => (x"9f",x"49",x"a2",x"d4"),
   727 => (x"c0",x"4c",x"49",x"69"),
   728 => (x"d0",x"9c",x"ff",x"ff"),
   729 => (x"c0",x"87",x"c2",x"34"),
   730 => (x"b3",x"49",x"74",x"4c"),
   731 => (x"ed",x"fd",x"49",x"73"),
   732 => (x"87",x"d9",x"ee",x"87"),
   733 => (x"5c",x"5b",x"5e",x"0e"),
   734 => (x"86",x"f4",x"0e",x"5d"),
   735 => (x"7e",x"c0",x"4a",x"71"),
   736 => (x"d8",x"02",x"9a",x"72"),
   737 => (x"e2",x"e5",x"c2",x"87"),
   738 => (x"c2",x"78",x"c0",x"48"),
   739 => (x"c2",x"48",x"da",x"e5"),
   740 => (x"78",x"bf",x"d3",x"f2"),
   741 => (x"48",x"de",x"e5",x"c2"),
   742 => (x"bf",x"cf",x"f2",x"c2"),
   743 => (x"c3",x"ee",x"c2",x"78"),
   744 => (x"c2",x"50",x"c0",x"48"),
   745 => (x"49",x"bf",x"f2",x"ed"),
   746 => (x"bf",x"e2",x"e5",x"c2"),
   747 => (x"03",x"aa",x"71",x"4a"),
   748 => (x"72",x"87",x"ca",x"c4"),
   749 => (x"05",x"99",x"cf",x"49"),
   750 => (x"c0",x"87",x"ea",x"c0"),
   751 => (x"c2",x"48",x"d0",x"f5"),
   752 => (x"78",x"bf",x"da",x"e5"),
   753 => (x"1e",x"e6",x"e5",x"c2"),
   754 => (x"bf",x"da",x"e5",x"c2"),
   755 => (x"da",x"e5",x"c2",x"49"),
   756 => (x"78",x"a1",x"c1",x"48"),
   757 => (x"f4",x"de",x"ff",x"71"),
   758 => (x"c0",x"86",x"c4",x"87"),
   759 => (x"c2",x"48",x"cc",x"f5"),
   760 => (x"cc",x"78",x"e6",x"e5"),
   761 => (x"cc",x"f5",x"c0",x"87"),
   762 => (x"e0",x"c0",x"48",x"bf"),
   763 => (x"d0",x"f5",x"c0",x"80"),
   764 => (x"e2",x"e5",x"c2",x"58"),
   765 => (x"80",x"c1",x"48",x"bf"),
   766 => (x"58",x"e6",x"e5",x"c2"),
   767 => (x"00",x"0d",x"4c",x"27"),
   768 => (x"bf",x"97",x"bf",x"00"),
   769 => (x"c2",x"02",x"9d",x"4d"),
   770 => (x"e5",x"c3",x"87",x"e3"),
   771 => (x"dc",x"c2",x"02",x"ad"),
   772 => (x"cc",x"f5",x"c0",x"87"),
   773 => (x"a3",x"cb",x"4b",x"bf"),
   774 => (x"cf",x"4c",x"11",x"49"),
   775 => (x"d2",x"c1",x"05",x"ac"),
   776 => (x"df",x"49",x"75",x"87"),
   777 => (x"cd",x"89",x"c1",x"99"),
   778 => (x"f6",x"ed",x"c2",x"91"),
   779 => (x"4a",x"a3",x"c1",x"81"),
   780 => (x"a3",x"c3",x"51",x"12"),
   781 => (x"c5",x"51",x"12",x"4a"),
   782 => (x"51",x"12",x"4a",x"a3"),
   783 => (x"12",x"4a",x"a3",x"c7"),
   784 => (x"4a",x"a3",x"c9",x"51"),
   785 => (x"a3",x"ce",x"51",x"12"),
   786 => (x"d0",x"51",x"12",x"4a"),
   787 => (x"51",x"12",x"4a",x"a3"),
   788 => (x"12",x"4a",x"a3",x"d2"),
   789 => (x"4a",x"a3",x"d4",x"51"),
   790 => (x"a3",x"d6",x"51",x"12"),
   791 => (x"d8",x"51",x"12",x"4a"),
   792 => (x"51",x"12",x"4a",x"a3"),
   793 => (x"12",x"4a",x"a3",x"dc"),
   794 => (x"4a",x"a3",x"de",x"51"),
   795 => (x"7e",x"c1",x"51",x"12"),
   796 => (x"74",x"87",x"fa",x"c0"),
   797 => (x"05",x"99",x"c8",x"49"),
   798 => (x"74",x"87",x"eb",x"c0"),
   799 => (x"05",x"99",x"d0",x"49"),
   800 => (x"66",x"dc",x"87",x"d1"),
   801 => (x"87",x"cb",x"c0",x"02"),
   802 => (x"66",x"dc",x"49",x"73"),
   803 => (x"02",x"98",x"70",x"0f"),
   804 => (x"6e",x"87",x"d3",x"c0"),
   805 => (x"87",x"c6",x"c0",x"05"),
   806 => (x"48",x"f6",x"ed",x"c2"),
   807 => (x"f5",x"c0",x"50",x"c0"),
   808 => (x"c2",x"48",x"bf",x"cc"),
   809 => (x"ee",x"c2",x"87",x"e1"),
   810 => (x"50",x"c0",x"48",x"c3"),
   811 => (x"f2",x"ed",x"c2",x"7e"),
   812 => (x"e5",x"c2",x"49",x"bf"),
   813 => (x"71",x"4a",x"bf",x"e2"),
   814 => (x"f6",x"fb",x"04",x"aa"),
   815 => (x"d3",x"f2",x"c2",x"87"),
   816 => (x"c8",x"c0",x"05",x"bf"),
   817 => (x"ee",x"ed",x"c2",x"87"),
   818 => (x"f8",x"c1",x"02",x"bf"),
   819 => (x"de",x"e5",x"c2",x"87"),
   820 => (x"fe",x"e8",x"49",x"bf"),
   821 => (x"c2",x"49",x"70",x"87"),
   822 => (x"c4",x"59",x"e2",x"e5"),
   823 => (x"e5",x"c2",x"48",x"a6"),
   824 => (x"c2",x"78",x"bf",x"de"),
   825 => (x"02",x"bf",x"ee",x"ed"),
   826 => (x"c4",x"87",x"d8",x"c0"),
   827 => (x"ff",x"cf",x"49",x"66"),
   828 => (x"99",x"f8",x"ff",x"ff"),
   829 => (x"c5",x"c0",x"02",x"a9"),
   830 => (x"c0",x"4c",x"c0",x"87"),
   831 => (x"4c",x"c1",x"87",x"e1"),
   832 => (x"c4",x"87",x"dc",x"c0"),
   833 => (x"ff",x"cf",x"49",x"66"),
   834 => (x"02",x"a9",x"99",x"f8"),
   835 => (x"c8",x"87",x"c8",x"c0"),
   836 => (x"78",x"c0",x"48",x"a6"),
   837 => (x"c8",x"87",x"c5",x"c0"),
   838 => (x"78",x"c1",x"48",x"a6"),
   839 => (x"74",x"4c",x"66",x"c8"),
   840 => (x"e0",x"c0",x"05",x"9c"),
   841 => (x"49",x"66",x"c4",x"87"),
   842 => (x"ed",x"c2",x"89",x"c2"),
   843 => (x"91",x"4a",x"bf",x"e6"),
   844 => (x"bf",x"ff",x"f1",x"c2"),
   845 => (x"da",x"e5",x"c2",x"4a"),
   846 => (x"78",x"a1",x"72",x"48"),
   847 => (x"48",x"e2",x"e5",x"c2"),
   848 => (x"de",x"f9",x"78",x"c0"),
   849 => (x"f4",x"48",x"c0",x"87"),
   850 => (x"87",x"ff",x"e6",x"8e"),
   851 => (x"00",x"00",x"00",x"00"),
   852 => (x"ff",x"ff",x"ff",x"ff"),
   853 => (x"00",x"00",x"0d",x"5c"),
   854 => (x"00",x"00",x"0d",x"65"),
   855 => (x"33",x"54",x"41",x"46"),
   856 => (x"20",x"20",x"20",x"32"),
   857 => (x"54",x"41",x"46",x"00"),
   858 => (x"20",x"20",x"36",x"31"),
   859 => (x"c2",x"1e",x"00",x"20"),
   860 => (x"48",x"bf",x"d8",x"f2"),
   861 => (x"c9",x"05",x"a8",x"dd"),
   862 => (x"e1",x"c2",x"c1",x"87"),
   863 => (x"4a",x"49",x"70",x"87"),
   864 => (x"d4",x"ff",x"87",x"c8"),
   865 => (x"78",x"ff",x"c3",x"48"),
   866 => (x"48",x"72",x"4a",x"68"),
   867 => (x"c2",x"1e",x"4f",x"26"),
   868 => (x"48",x"bf",x"d8",x"f2"),
   869 => (x"c6",x"05",x"a8",x"dd"),
   870 => (x"ed",x"c1",x"c1",x"87"),
   871 => (x"ff",x"87",x"d9",x"87"),
   872 => (x"ff",x"c3",x"48",x"d4"),
   873 => (x"48",x"d0",x"ff",x"78"),
   874 => (x"ff",x"78",x"e1",x"c0"),
   875 => (x"78",x"d4",x"48",x"d4"),
   876 => (x"48",x"d7",x"f2",x"c2"),
   877 => (x"50",x"bf",x"d4",x"ff"),
   878 => (x"ff",x"1e",x"4f",x"26"),
   879 => (x"e0",x"c0",x"48",x"d0"),
   880 => (x"1e",x"4f",x"26",x"78"),
   881 => (x"70",x"87",x"e7",x"fe"),
   882 => (x"c6",x"02",x"99",x"49"),
   883 => (x"a9",x"fb",x"c0",x"87"),
   884 => (x"71",x"87",x"f1",x"05"),
   885 => (x"0e",x"4f",x"26",x"48"),
   886 => (x"0e",x"5c",x"5b",x"5e"),
   887 => (x"4c",x"c0",x"4b",x"71"),
   888 => (x"70",x"87",x"cb",x"fe"),
   889 => (x"c0",x"02",x"99",x"49"),
   890 => (x"ec",x"c0",x"87",x"f9"),
   891 => (x"f2",x"c0",x"02",x"a9"),
   892 => (x"a9",x"fb",x"c0",x"87"),
   893 => (x"87",x"eb",x"c0",x"02"),
   894 => (x"ac",x"b7",x"66",x"cc"),
   895 => (x"d0",x"87",x"c7",x"03"),
   896 => (x"87",x"c2",x"02",x"66"),
   897 => (x"99",x"71",x"53",x"71"),
   898 => (x"c1",x"87",x"c2",x"02"),
   899 => (x"87",x"de",x"fd",x"84"),
   900 => (x"02",x"99",x"49",x"70"),
   901 => (x"ec",x"c0",x"87",x"cd"),
   902 => (x"87",x"c7",x"02",x"a9"),
   903 => (x"05",x"a9",x"fb",x"c0"),
   904 => (x"d0",x"87",x"d5",x"ff"),
   905 => (x"87",x"c3",x"02",x"66"),
   906 => (x"c0",x"7b",x"97",x"c0"),
   907 => (x"c4",x"05",x"a9",x"ec"),
   908 => (x"c5",x"4a",x"74",x"87"),
   909 => (x"c0",x"4a",x"74",x"87"),
   910 => (x"48",x"72",x"8a",x"0a"),
   911 => (x"4d",x"26",x"87",x"c2"),
   912 => (x"4b",x"26",x"4c",x"26"),
   913 => (x"fc",x"1e",x"4f",x"26"),
   914 => (x"49",x"70",x"87",x"e4"),
   915 => (x"aa",x"f0",x"c0",x"4a"),
   916 => (x"c0",x"87",x"c9",x"04"),
   917 => (x"c3",x"01",x"aa",x"f9"),
   918 => (x"8a",x"f0",x"c0",x"87"),
   919 => (x"04",x"aa",x"c1",x"c1"),
   920 => (x"da",x"c1",x"87",x"c9"),
   921 => (x"87",x"c3",x"01",x"aa"),
   922 => (x"72",x"8a",x"f7",x"c0"),
   923 => (x"0e",x"4f",x"26",x"48"),
   924 => (x"0e",x"5c",x"5b",x"5e"),
   925 => (x"d4",x"ff",x"4a",x"71"),
   926 => (x"c0",x"49",x"72",x"4c"),
   927 => (x"4b",x"70",x"87",x"e9"),
   928 => (x"87",x"c2",x"02",x"9b"),
   929 => (x"d0",x"ff",x"8b",x"c1"),
   930 => (x"c1",x"78",x"c5",x"48"),
   931 => (x"49",x"73",x"7c",x"d5"),
   932 => (x"e7",x"c1",x"31",x"c6"),
   933 => (x"4a",x"bf",x"97",x"d0"),
   934 => (x"70",x"b0",x"71",x"48"),
   935 => (x"48",x"d0",x"ff",x"7c"),
   936 => (x"48",x"73",x"78",x"c4"),
   937 => (x"0e",x"87",x"d9",x"fe"),
   938 => (x"5d",x"5c",x"5b",x"5e"),
   939 => (x"71",x"86",x"f8",x"0e"),
   940 => (x"c0",x"7e",x"c0",x"4b"),
   941 => (x"bf",x"97",x"cd",x"fe"),
   942 => (x"c0",x"05",x"99",x"49"),
   943 => (x"a3",x"c8",x"87",x"ee"),
   944 => (x"49",x"69",x"97",x"49"),
   945 => (x"05",x"a9",x"c1",x"c1"),
   946 => (x"a3",x"c9",x"87",x"dd"),
   947 => (x"49",x"69",x"97",x"49"),
   948 => (x"05",x"a9",x"d2",x"c1"),
   949 => (x"a3",x"ca",x"87",x"d1"),
   950 => (x"49",x"69",x"97",x"49"),
   951 => (x"05",x"a9",x"c3",x"c1"),
   952 => (x"48",x"df",x"87",x"c5"),
   953 => (x"c0",x"87",x"e1",x"c2"),
   954 => (x"87",x"dc",x"c2",x"48"),
   955 => (x"c0",x"87",x"df",x"fa"),
   956 => (x"cd",x"fe",x"c0",x"4c"),
   957 => (x"c0",x"49",x"bf",x"97"),
   958 => (x"87",x"cf",x"04",x"a9"),
   959 => (x"c1",x"87",x"c4",x"fb"),
   960 => (x"cd",x"fe",x"c0",x"84"),
   961 => (x"ac",x"49",x"bf",x"97"),
   962 => (x"c0",x"87",x"f1",x"06"),
   963 => (x"bf",x"97",x"cd",x"fe"),
   964 => (x"f9",x"87",x"cf",x"02"),
   965 => (x"49",x"70",x"87",x"d8"),
   966 => (x"87",x"c6",x"02",x"99"),
   967 => (x"05",x"a9",x"ec",x"c0"),
   968 => (x"4c",x"c0",x"87",x"f1"),
   969 => (x"70",x"87",x"c7",x"f9"),
   970 => (x"87",x"c2",x"f9",x"4d"),
   971 => (x"f8",x"58",x"a6",x"c8"),
   972 => (x"4a",x"70",x"87",x"fc"),
   973 => (x"a3",x"c8",x"84",x"c1"),
   974 => (x"49",x"69",x"97",x"49"),
   975 => (x"87",x"c7",x"02",x"ad"),
   976 => (x"05",x"ad",x"ff",x"c0"),
   977 => (x"c9",x"87",x"e7",x"c0"),
   978 => (x"69",x"97",x"49",x"a3"),
   979 => (x"a9",x"66",x"c4",x"49"),
   980 => (x"48",x"87",x"c7",x"02"),
   981 => (x"05",x"a8",x"ff",x"c0"),
   982 => (x"a3",x"ca",x"87",x"d4"),
   983 => (x"49",x"69",x"97",x"49"),
   984 => (x"87",x"c6",x"02",x"aa"),
   985 => (x"05",x"aa",x"ff",x"c0"),
   986 => (x"7e",x"c1",x"87",x"c4"),
   987 => (x"ec",x"c0",x"87",x"d0"),
   988 => (x"87",x"c6",x"02",x"ad"),
   989 => (x"05",x"ad",x"fb",x"c0"),
   990 => (x"4c",x"c0",x"87",x"c4"),
   991 => (x"02",x"6e",x"7e",x"c1"),
   992 => (x"f8",x"87",x"e1",x"fe"),
   993 => (x"48",x"74",x"87",x"f4"),
   994 => (x"f1",x"fa",x"8e",x"f8"),
   995 => (x"5e",x"0e",x"00",x"87"),
   996 => (x"0e",x"5d",x"5c",x"5b"),
   997 => (x"4d",x"71",x"86",x"f8"),
   998 => (x"75",x"4b",x"d4",x"ff"),
   999 => (x"dc",x"f2",x"c2",x"1e"),
  1000 => (x"e0",x"df",x"ff",x"49"),
  1001 => (x"70",x"86",x"c4",x"87"),
  1002 => (x"fb",x"c4",x"02",x"98"),
  1003 => (x"d2",x"e7",x"c1",x"87"),
  1004 => (x"49",x"75",x"7e",x"bf"),
  1005 => (x"de",x"87",x"f8",x"fa"),
  1006 => (x"eb",x"c0",x"05",x"a8"),
  1007 => (x"c0",x"49",x"75",x"87"),
  1008 => (x"70",x"87",x"f9",x"f6"),
  1009 => (x"87",x"db",x"02",x"98"),
  1010 => (x"bf",x"c0",x"f7",x"c2"),
  1011 => (x"49",x"e1",x"c0",x"1e"),
  1012 => (x"87",x"c8",x"f4",x"c0"),
  1013 => (x"e7",x"c1",x"86",x"c4"),
  1014 => (x"50",x"c0",x"48",x"d0"),
  1015 => (x"49",x"cc",x"f7",x"c2"),
  1016 => (x"c1",x"87",x"eb",x"fe"),
  1017 => (x"87",x"c2",x"c4",x"48"),
  1018 => (x"c5",x"48",x"d0",x"ff"),
  1019 => (x"7b",x"d6",x"c1",x"78"),
  1020 => (x"a2",x"75",x"4a",x"c0"),
  1021 => (x"c1",x"7b",x"11",x"49"),
  1022 => (x"aa",x"b7",x"cb",x"82"),
  1023 => (x"cc",x"87",x"f3",x"04"),
  1024 => (x"7b",x"ff",x"c3",x"4a"),
  1025 => (x"e0",x"c0",x"82",x"c1"),
  1026 => (x"f4",x"04",x"aa",x"b7"),
  1027 => (x"48",x"d0",x"ff",x"87"),
  1028 => (x"ff",x"c3",x"78",x"c4"),
  1029 => (x"c1",x"78",x"c5",x"7b"),
  1030 => (x"7b",x"c1",x"7b",x"d3"),
  1031 => (x"48",x"6e",x"78",x"c4"),
  1032 => (x"06",x"a8",x"b7",x"c0"),
  1033 => (x"c2",x"87",x"f0",x"c2"),
  1034 => (x"4c",x"bf",x"e4",x"f2"),
  1035 => (x"88",x"74",x"48",x"6e"),
  1036 => (x"9c",x"74",x"7e",x"70"),
  1037 => (x"87",x"fd",x"c1",x"02"),
  1038 => (x"4d",x"e6",x"e5",x"c2"),
  1039 => (x"c8",x"48",x"a6",x"c4"),
  1040 => (x"c0",x"8c",x"78",x"c0"),
  1041 => (x"c6",x"03",x"ac",x"b7"),
  1042 => (x"a4",x"c0",x"c8",x"87"),
  1043 => (x"c2",x"4c",x"c0",x"78"),
  1044 => (x"bf",x"97",x"d7",x"f2"),
  1045 => (x"02",x"99",x"d0",x"49"),
  1046 => (x"1e",x"c0",x"87",x"d1"),
  1047 => (x"49",x"dc",x"f2",x"c2"),
  1048 => (x"c4",x"87",x"d5",x"e1"),
  1049 => (x"4a",x"49",x"70",x"86"),
  1050 => (x"c2",x"87",x"ee",x"c0"),
  1051 => (x"c2",x"1e",x"e6",x"e5"),
  1052 => (x"e1",x"49",x"dc",x"f2"),
  1053 => (x"86",x"c4",x"87",x"c2"),
  1054 => (x"ff",x"4a",x"49",x"70"),
  1055 => (x"c5",x"c8",x"48",x"d0"),
  1056 => (x"7b",x"d4",x"c1",x"78"),
  1057 => (x"66",x"c4",x"7b",x"15"),
  1058 => (x"c8",x"88",x"c1",x"48"),
  1059 => (x"98",x"70",x"58",x"a6"),
  1060 => (x"87",x"f0",x"ff",x"05"),
  1061 => (x"c4",x"48",x"d0",x"ff"),
  1062 => (x"05",x"9a",x"72",x"78"),
  1063 => (x"48",x"c0",x"87",x"c5"),
  1064 => (x"c1",x"87",x"c7",x"c1"),
  1065 => (x"dc",x"f2",x"c2",x"1e"),
  1066 => (x"f1",x"de",x"ff",x"49"),
  1067 => (x"74",x"86",x"c4",x"87"),
  1068 => (x"c3",x"fe",x"05",x"9c"),
  1069 => (x"c0",x"48",x"6e",x"87"),
  1070 => (x"d1",x"06",x"a8",x"b7"),
  1071 => (x"dc",x"f2",x"c2",x"87"),
  1072 => (x"d0",x"78",x"c0",x"48"),
  1073 => (x"f4",x"78",x"c0",x"80"),
  1074 => (x"e8",x"f2",x"c2",x"80"),
  1075 => (x"48",x"6e",x"78",x"bf"),
  1076 => (x"01",x"a8",x"b7",x"c0"),
  1077 => (x"ff",x"87",x"d0",x"fd"),
  1078 => (x"78",x"c5",x"48",x"d0"),
  1079 => (x"c0",x"7b",x"d3",x"c1"),
  1080 => (x"c1",x"78",x"c4",x"7b"),
  1081 => (x"87",x"c2",x"c0",x"48"),
  1082 => (x"8e",x"f8",x"48",x"c0"),
  1083 => (x"4c",x"26",x"4d",x"26"),
  1084 => (x"4f",x"26",x"4b",x"26"),
  1085 => (x"5c",x"5b",x"5e",x"0e"),
  1086 => (x"71",x"1e",x"0e",x"5d"),
  1087 => (x"4d",x"4c",x"c0",x"4b"),
  1088 => (x"e8",x"c0",x"04",x"ab"),
  1089 => (x"e7",x"fa",x"c0",x"87"),
  1090 => (x"02",x"9d",x"75",x"1e"),
  1091 => (x"4a",x"c0",x"87",x"c4"),
  1092 => (x"4a",x"c1",x"87",x"c2"),
  1093 => (x"db",x"e9",x"49",x"72"),
  1094 => (x"70",x"86",x"c4",x"87"),
  1095 => (x"6e",x"84",x"c1",x"7e"),
  1096 => (x"73",x"87",x"c2",x"05"),
  1097 => (x"73",x"85",x"c1",x"4c"),
  1098 => (x"d8",x"ff",x"06",x"ac"),
  1099 => (x"26",x"48",x"6e",x"87"),
  1100 => (x"1e",x"87",x"f9",x"fe"),
  1101 => (x"66",x"c4",x"4a",x"71"),
  1102 => (x"72",x"87",x"c5",x"05"),
  1103 => (x"87",x"ce",x"f9",x"49"),
  1104 => (x"5e",x"0e",x"4f",x"26"),
  1105 => (x"0e",x"5d",x"5c",x"5b"),
  1106 => (x"49",x"4c",x"71",x"1e"),
  1107 => (x"f3",x"c2",x"91",x"de"),
  1108 => (x"85",x"71",x"4d",x"c4"),
  1109 => (x"c1",x"02",x"6d",x"97"),
  1110 => (x"f2",x"c2",x"87",x"dc"),
  1111 => (x"74",x"4a",x"bf",x"f0"),
  1112 => (x"fe",x"49",x"72",x"82"),
  1113 => (x"7e",x"70",x"87",x"ce"),
  1114 => (x"f2",x"c0",x"02",x"6e"),
  1115 => (x"f8",x"f2",x"c2",x"87"),
  1116 => (x"cb",x"4a",x"6e",x"4b"),
  1117 => (x"ef",x"fc",x"fe",x"49"),
  1118 => (x"cb",x"4b",x"74",x"87"),
  1119 => (x"e4",x"e7",x"c1",x"93"),
  1120 => (x"c1",x"83",x"c4",x"83"),
  1121 => (x"74",x"7b",x"fa",x"c6"),
  1122 => (x"d0",x"cb",x"c1",x"49"),
  1123 => (x"c1",x"7b",x"75",x"87"),
  1124 => (x"bf",x"97",x"d1",x"e7"),
  1125 => (x"f2",x"c2",x"1e",x"49"),
  1126 => (x"d6",x"fe",x"49",x"f8"),
  1127 => (x"74",x"86",x"c4",x"87"),
  1128 => (x"f8",x"ca",x"c1",x"49"),
  1129 => (x"c1",x"49",x"c0",x"87"),
  1130 => (x"c2",x"87",x"d7",x"cc"),
  1131 => (x"c0",x"48",x"d8",x"f2"),
  1132 => (x"dd",x"49",x"c1",x"78"),
  1133 => (x"fc",x"26",x"87",x"d9"),
  1134 => (x"6f",x"4c",x"87",x"f2"),
  1135 => (x"6e",x"69",x"64",x"61"),
  1136 => (x"2e",x"2e",x"2e",x"67"),
  1137 => (x"5b",x"5e",x"0e",x"00"),
  1138 => (x"4b",x"71",x"0e",x"5c"),
  1139 => (x"f0",x"f2",x"c2",x"4a"),
  1140 => (x"49",x"72",x"82",x"bf"),
  1141 => (x"70",x"87",x"dd",x"fc"),
  1142 => (x"c4",x"02",x"9c",x"4c"),
  1143 => (x"db",x"e5",x"49",x"87"),
  1144 => (x"f0",x"f2",x"c2",x"87"),
  1145 => (x"c1",x"78",x"c0",x"48"),
  1146 => (x"87",x"e3",x"dc",x"49"),
  1147 => (x"0e",x"87",x"ff",x"fb"),
  1148 => (x"5d",x"5c",x"5b",x"5e"),
  1149 => (x"c2",x"86",x"f4",x"0e"),
  1150 => (x"c0",x"4d",x"e6",x"e5"),
  1151 => (x"48",x"a6",x"c4",x"4c"),
  1152 => (x"f2",x"c2",x"78",x"c0"),
  1153 => (x"c0",x"49",x"bf",x"f0"),
  1154 => (x"c1",x"c1",x"06",x"a9"),
  1155 => (x"e6",x"e5",x"c2",x"87"),
  1156 => (x"c0",x"02",x"98",x"48"),
  1157 => (x"fa",x"c0",x"87",x"f8"),
  1158 => (x"66",x"c8",x"1e",x"e7"),
  1159 => (x"c4",x"87",x"c7",x"02"),
  1160 => (x"78",x"c0",x"48",x"a6"),
  1161 => (x"a6",x"c4",x"87",x"c5"),
  1162 => (x"c4",x"78",x"c1",x"48"),
  1163 => (x"c3",x"e5",x"49",x"66"),
  1164 => (x"70",x"86",x"c4",x"87"),
  1165 => (x"c4",x"84",x"c1",x"4d"),
  1166 => (x"80",x"c1",x"48",x"66"),
  1167 => (x"c2",x"58",x"a6",x"c8"),
  1168 => (x"49",x"bf",x"f0",x"f2"),
  1169 => (x"87",x"c6",x"03",x"ac"),
  1170 => (x"ff",x"05",x"9d",x"75"),
  1171 => (x"4c",x"c0",x"87",x"c8"),
  1172 => (x"c3",x"02",x"9d",x"75"),
  1173 => (x"fa",x"c0",x"87",x"e0"),
  1174 => (x"66",x"c8",x"1e",x"e7"),
  1175 => (x"cc",x"87",x"c7",x"02"),
  1176 => (x"78",x"c0",x"48",x"a6"),
  1177 => (x"a6",x"cc",x"87",x"c5"),
  1178 => (x"cc",x"78",x"c1",x"48"),
  1179 => (x"c3",x"e4",x"49",x"66"),
  1180 => (x"70",x"86",x"c4",x"87"),
  1181 => (x"c2",x"02",x"6e",x"7e"),
  1182 => (x"49",x"6e",x"87",x"e9"),
  1183 => (x"69",x"97",x"81",x"cb"),
  1184 => (x"02",x"99",x"d0",x"49"),
  1185 => (x"c1",x"87",x"d6",x"c1"),
  1186 => (x"74",x"4a",x"c5",x"c7"),
  1187 => (x"c1",x"91",x"cb",x"49"),
  1188 => (x"72",x"81",x"e4",x"e7"),
  1189 => (x"c3",x"81",x"c8",x"79"),
  1190 => (x"49",x"74",x"51",x"ff"),
  1191 => (x"f3",x"c2",x"91",x"de"),
  1192 => (x"85",x"71",x"4d",x"c4"),
  1193 => (x"7d",x"97",x"c1",x"c2"),
  1194 => (x"c0",x"49",x"a5",x"c1"),
  1195 => (x"ed",x"c2",x"51",x"e0"),
  1196 => (x"02",x"bf",x"97",x"f6"),
  1197 => (x"84",x"c1",x"87",x"d2"),
  1198 => (x"c2",x"4b",x"a5",x"c2"),
  1199 => (x"db",x"4a",x"f6",x"ed"),
  1200 => (x"e3",x"f7",x"fe",x"49"),
  1201 => (x"87",x"db",x"c1",x"87"),
  1202 => (x"c0",x"49",x"a5",x"cd"),
  1203 => (x"c2",x"84",x"c1",x"51"),
  1204 => (x"4a",x"6e",x"4b",x"a5"),
  1205 => (x"f7",x"fe",x"49",x"cb"),
  1206 => (x"c6",x"c1",x"87",x"ce"),
  1207 => (x"c2",x"c5",x"c1",x"87"),
  1208 => (x"cb",x"49",x"74",x"4a"),
  1209 => (x"e4",x"e7",x"c1",x"91"),
  1210 => (x"c2",x"79",x"72",x"81"),
  1211 => (x"bf",x"97",x"f6",x"ed"),
  1212 => (x"74",x"87",x"d8",x"02"),
  1213 => (x"c1",x"91",x"de",x"49"),
  1214 => (x"c4",x"f3",x"c2",x"84"),
  1215 => (x"c2",x"83",x"71",x"4b"),
  1216 => (x"dd",x"4a",x"f6",x"ed"),
  1217 => (x"df",x"f6",x"fe",x"49"),
  1218 => (x"74",x"87",x"d8",x"87"),
  1219 => (x"c2",x"93",x"de",x"4b"),
  1220 => (x"cb",x"83",x"c4",x"f3"),
  1221 => (x"51",x"c0",x"49",x"a3"),
  1222 => (x"6e",x"73",x"84",x"c1"),
  1223 => (x"fe",x"49",x"cb",x"4a"),
  1224 => (x"c4",x"87",x"c5",x"f6"),
  1225 => (x"80",x"c1",x"48",x"66"),
  1226 => (x"c7",x"58",x"a6",x"c8"),
  1227 => (x"c5",x"c0",x"03",x"ac"),
  1228 => (x"fc",x"05",x"6e",x"87"),
  1229 => (x"48",x"74",x"87",x"e0"),
  1230 => (x"ef",x"f6",x"8e",x"f4"),
  1231 => (x"1e",x"73",x"1e",x"87"),
  1232 => (x"cb",x"49",x"4b",x"71"),
  1233 => (x"e4",x"e7",x"c1",x"91"),
  1234 => (x"4a",x"a1",x"c8",x"81"),
  1235 => (x"48",x"d0",x"e7",x"c1"),
  1236 => (x"a1",x"c9",x"50",x"12"),
  1237 => (x"cd",x"fe",x"c0",x"4a"),
  1238 => (x"ca",x"50",x"12",x"48"),
  1239 => (x"d1",x"e7",x"c1",x"81"),
  1240 => (x"c1",x"50",x"11",x"48"),
  1241 => (x"bf",x"97",x"d1",x"e7"),
  1242 => (x"49",x"c0",x"1e",x"49"),
  1243 => (x"c2",x"87",x"c4",x"f7"),
  1244 => (x"de",x"48",x"d8",x"f2"),
  1245 => (x"d6",x"49",x"c1",x"78"),
  1246 => (x"f5",x"26",x"87",x"d5"),
  1247 => (x"71",x"1e",x"87",x"f2"),
  1248 => (x"91",x"cb",x"49",x"4a"),
  1249 => (x"81",x"e4",x"e7",x"c1"),
  1250 => (x"48",x"11",x"81",x"c8"),
  1251 => (x"58",x"dc",x"f2",x"c2"),
  1252 => (x"48",x"f0",x"f2",x"c2"),
  1253 => (x"49",x"c1",x"78",x"c0"),
  1254 => (x"26",x"87",x"f4",x"d5"),
  1255 => (x"49",x"c0",x"1e",x"4f"),
  1256 => (x"87",x"de",x"c4",x"c1"),
  1257 => (x"71",x"1e",x"4f",x"26"),
  1258 => (x"87",x"d2",x"02",x"99"),
  1259 => (x"48",x"f9",x"e8",x"c1"),
  1260 => (x"80",x"f7",x"50",x"c0"),
  1261 => (x"40",x"fe",x"cd",x"c1"),
  1262 => (x"78",x"dd",x"e7",x"c1"),
  1263 => (x"e8",x"c1",x"87",x"ce"),
  1264 => (x"e7",x"c1",x"48",x"f5"),
  1265 => (x"80",x"fc",x"78",x"d6"),
  1266 => (x"78",x"dd",x"ce",x"c1"),
  1267 => (x"5e",x"0e",x"4f",x"26"),
  1268 => (x"71",x"0e",x"5c",x"5b"),
  1269 => (x"92",x"cb",x"4a",x"4c"),
  1270 => (x"82",x"e4",x"e7",x"c1"),
  1271 => (x"c9",x"49",x"a2",x"c8"),
  1272 => (x"6b",x"97",x"4b",x"a2"),
  1273 => (x"69",x"97",x"1e",x"4b"),
  1274 => (x"82",x"ca",x"1e",x"49"),
  1275 => (x"e5",x"c0",x"49",x"12"),
  1276 => (x"49",x"c0",x"87",x"ca"),
  1277 => (x"74",x"87",x"d8",x"d4"),
  1278 => (x"e0",x"c1",x"c1",x"49"),
  1279 => (x"f3",x"8e",x"f8",x"87"),
  1280 => (x"73",x"1e",x"87",x"ec"),
  1281 => (x"49",x"4b",x"71",x"1e"),
  1282 => (x"73",x"87",x"c3",x"ff"),
  1283 => (x"87",x"fe",x"fe",x"49"),
  1284 => (x"1e",x"87",x"dd",x"f3"),
  1285 => (x"4b",x"71",x"1e",x"73"),
  1286 => (x"02",x"4a",x"a3",x"c6"),
  1287 => (x"8a",x"c1",x"87",x"db"),
  1288 => (x"8a",x"87",x"d6",x"02"),
  1289 => (x"87",x"da",x"c1",x"02"),
  1290 => (x"fc",x"c0",x"02",x"8a"),
  1291 => (x"c0",x"02",x"8a",x"87"),
  1292 => (x"02",x"8a",x"87",x"e1"),
  1293 => (x"db",x"c1",x"87",x"cb"),
  1294 => (x"fd",x"49",x"c7",x"87"),
  1295 => (x"de",x"c1",x"87",x"c0"),
  1296 => (x"f0",x"f2",x"c2",x"87"),
  1297 => (x"cb",x"c1",x"02",x"bf"),
  1298 => (x"88",x"c1",x"48",x"87"),
  1299 => (x"58",x"f4",x"f2",x"c2"),
  1300 => (x"c2",x"87",x"c1",x"c1"),
  1301 => (x"02",x"bf",x"f4",x"f2"),
  1302 => (x"c2",x"87",x"f9",x"c0"),
  1303 => (x"48",x"bf",x"f0",x"f2"),
  1304 => (x"f2",x"c2",x"80",x"c1"),
  1305 => (x"eb",x"c0",x"58",x"f4"),
  1306 => (x"f0",x"f2",x"c2",x"87"),
  1307 => (x"89",x"c6",x"49",x"bf"),
  1308 => (x"59",x"f4",x"f2",x"c2"),
  1309 => (x"03",x"a9",x"b7",x"c0"),
  1310 => (x"f2",x"c2",x"87",x"da"),
  1311 => (x"78",x"c0",x"48",x"f0"),
  1312 => (x"f2",x"c2",x"87",x"d2"),
  1313 => (x"cb",x"02",x"bf",x"f4"),
  1314 => (x"f0",x"f2",x"c2",x"87"),
  1315 => (x"80",x"c6",x"48",x"bf"),
  1316 => (x"58",x"f4",x"f2",x"c2"),
  1317 => (x"f6",x"d1",x"49",x"c0"),
  1318 => (x"c0",x"49",x"73",x"87"),
  1319 => (x"f1",x"87",x"fe",x"fe"),
  1320 => (x"73",x"1e",x"87",x"ce"),
  1321 => (x"c2",x"4b",x"71",x"1e"),
  1322 => (x"dd",x"48",x"d8",x"f2"),
  1323 => (x"d1",x"49",x"c0",x"78"),
  1324 => (x"49",x"73",x"87",x"dd"),
  1325 => (x"87",x"e5",x"fe",x"c0"),
  1326 => (x"0e",x"87",x"f5",x"f0"),
  1327 => (x"5d",x"5c",x"5b",x"5e"),
  1328 => (x"86",x"cc",x"ff",x"0e"),
  1329 => (x"c8",x"59",x"a6",x"d8"),
  1330 => (x"78",x"c0",x"48",x"a6"),
  1331 => (x"c8",x"c1",x"80",x"c4"),
  1332 => (x"80",x"c4",x"78",x"66"),
  1333 => (x"f2",x"c2",x"78",x"c1"),
  1334 => (x"78",x"c1",x"48",x"f4"),
  1335 => (x"bf",x"d8",x"f2",x"c2"),
  1336 => (x"05",x"a8",x"de",x"48"),
  1337 => (x"c6",x"f4",x"87",x"cb"),
  1338 => (x"cc",x"49",x"70",x"87"),
  1339 => (x"d0",x"cf",x"59",x"a6"),
  1340 => (x"87",x"da",x"e2",x"87"),
  1341 => (x"e1",x"87",x"cc",x"e3"),
  1342 => (x"4c",x"70",x"87",x"f4"),
  1343 => (x"c1",x"05",x"66",x"d4"),
  1344 => (x"c4",x"c1",x"87",x"fc"),
  1345 => (x"80",x"c4",x"48",x"66"),
  1346 => (x"a6",x"c4",x"7e",x"70"),
  1347 => (x"78",x"bf",x"6e",x"48"),
  1348 => (x"e3",x"c1",x"1e",x"72"),
  1349 => (x"66",x"c8",x"48",x"f6"),
  1350 => (x"4a",x"a1",x"c8",x"49"),
  1351 => (x"aa",x"71",x"41",x"20"),
  1352 => (x"10",x"87",x"f9",x"05"),
  1353 => (x"c1",x"4a",x"26",x"51"),
  1354 => (x"c1",x"48",x"66",x"c4"),
  1355 => (x"6e",x"78",x"fd",x"cc"),
  1356 => (x"81",x"c7",x"49",x"bf"),
  1357 => (x"c4",x"c1",x"51",x"74"),
  1358 => (x"81",x"c8",x"49",x"66"),
  1359 => (x"c4",x"c1",x"51",x"c1"),
  1360 => (x"81",x"c9",x"49",x"66"),
  1361 => (x"c4",x"c1",x"51",x"c0"),
  1362 => (x"81",x"ca",x"49",x"66"),
  1363 => (x"fb",x"c0",x"51",x"c0"),
  1364 => (x"87",x"cf",x"02",x"ac"),
  1365 => (x"1e",x"d8",x"1e",x"c1"),
  1366 => (x"49",x"bf",x"66",x"c8"),
  1367 => (x"f6",x"e1",x"81",x"c8"),
  1368 => (x"c1",x"86",x"c8",x"87"),
  1369 => (x"c0",x"48",x"66",x"c8"),
  1370 => (x"87",x"c7",x"01",x"a8"),
  1371 => (x"c1",x"48",x"a6",x"c8"),
  1372 => (x"c1",x"87",x"ce",x"78"),
  1373 => (x"c1",x"48",x"66",x"c8"),
  1374 => (x"58",x"a6",x"d0",x"88"),
  1375 => (x"c2",x"e1",x"87",x"c3"),
  1376 => (x"48",x"a6",x"d8",x"87"),
  1377 => (x"9c",x"74",x"78",x"c2"),
  1378 => (x"87",x"f1",x"cc",x"02"),
  1379 => (x"c1",x"48",x"66",x"c8"),
  1380 => (x"03",x"a8",x"66",x"cc"),
  1381 => (x"dc",x"87",x"e6",x"cc"),
  1382 => (x"78",x"c0",x"48",x"a6"),
  1383 => (x"78",x"c0",x"80",x"c4"),
  1384 => (x"87",x"ca",x"df",x"ff"),
  1385 => (x"66",x"d4",x"4c",x"70"),
  1386 => (x"05",x"a8",x"dd",x"48"),
  1387 => (x"e0",x"c0",x"87",x"c7"),
  1388 => (x"66",x"d4",x"48",x"a6"),
  1389 => (x"ac",x"d0",x"c1",x"78"),
  1390 => (x"87",x"eb",x"c0",x"05"),
  1391 => (x"87",x"ee",x"de",x"ff"),
  1392 => (x"87",x"ea",x"de",x"ff"),
  1393 => (x"ec",x"c0",x"4c",x"70"),
  1394 => (x"87",x"c6",x"05",x"ac"),
  1395 => (x"87",x"f3",x"df",x"ff"),
  1396 => (x"d0",x"c1",x"4c",x"70"),
  1397 => (x"87",x"c8",x"05",x"ac"),
  1398 => (x"c1",x"48",x"66",x"d0"),
  1399 => (x"58",x"a6",x"d4",x"80"),
  1400 => (x"02",x"ac",x"d0",x"c1"),
  1401 => (x"c0",x"87",x"d5",x"ff"),
  1402 => (x"d4",x"48",x"a6",x"e4"),
  1403 => (x"e0",x"c0",x"78",x"66"),
  1404 => (x"e4",x"c0",x"48",x"66"),
  1405 => (x"ca",x"05",x"a8",x"66"),
  1406 => (x"e8",x"c0",x"87",x"d5"),
  1407 => (x"78",x"c0",x"48",x"a6"),
  1408 => (x"c0",x"80",x"dc",x"ff"),
  1409 => (x"c0",x"4d",x"74",x"78"),
  1410 => (x"c9",x"02",x"8d",x"fb"),
  1411 => (x"8d",x"c9",x"87",x"db"),
  1412 => (x"c2",x"87",x"db",x"02"),
  1413 => (x"f7",x"c1",x"02",x"8d"),
  1414 => (x"02",x"8d",x"c9",x"87"),
  1415 => (x"c4",x"87",x"d8",x"c4"),
  1416 => (x"c1",x"c1",x"02",x"8d"),
  1417 => (x"02",x"8d",x"c1",x"87"),
  1418 => (x"c8",x"87",x"cc",x"c4"),
  1419 => (x"66",x"c8",x"87",x"f5"),
  1420 => (x"c1",x"91",x"cb",x"49"),
  1421 => (x"c4",x"81",x"66",x"c4"),
  1422 => (x"7e",x"6a",x"4a",x"a1"),
  1423 => (x"e4",x"c1",x"1e",x"71"),
  1424 => (x"66",x"c4",x"48",x"c2"),
  1425 => (x"4a",x"a1",x"cc",x"49"),
  1426 => (x"aa",x"71",x"41",x"20"),
  1427 => (x"87",x"f8",x"ff",x"05"),
  1428 => (x"49",x"26",x"51",x"10"),
  1429 => (x"79",x"e2",x"d2",x"c1"),
  1430 => (x"87",x"d2",x"dc",x"ff"),
  1431 => (x"a6",x"c4",x"4c",x"70"),
  1432 => (x"c8",x"78",x"c1",x"48"),
  1433 => (x"a6",x"dc",x"87",x"c3"),
  1434 => (x"78",x"f0",x"c0",x"48"),
  1435 => (x"87",x"fe",x"db",x"ff"),
  1436 => (x"ec",x"c0",x"4c",x"70"),
  1437 => (x"c4",x"c0",x"02",x"ac"),
  1438 => (x"a6",x"e0",x"c0",x"87"),
  1439 => (x"ac",x"ec",x"c0",x"5c"),
  1440 => (x"ff",x"87",x"cd",x"02"),
  1441 => (x"70",x"87",x"e7",x"db"),
  1442 => (x"ac",x"ec",x"c0",x"4c"),
  1443 => (x"87",x"f3",x"ff",x"05"),
  1444 => (x"02",x"ac",x"ec",x"c0"),
  1445 => (x"ff",x"87",x"c4",x"c0"),
  1446 => (x"c0",x"87",x"d3",x"db"),
  1447 => (x"d0",x"1e",x"ca",x"1e"),
  1448 => (x"91",x"cb",x"49",x"66"),
  1449 => (x"48",x"66",x"cc",x"c1"),
  1450 => (x"a6",x"cc",x"80",x"71"),
  1451 => (x"48",x"66",x"c8",x"58"),
  1452 => (x"a6",x"d0",x"80",x"c4"),
  1453 => (x"bf",x"66",x"cc",x"58"),
  1454 => (x"da",x"dc",x"ff",x"49"),
  1455 => (x"de",x"1e",x"c1",x"87"),
  1456 => (x"bf",x"66",x"d4",x"1e"),
  1457 => (x"ce",x"dc",x"ff",x"49"),
  1458 => (x"70",x"86",x"d0",x"87"),
  1459 => (x"89",x"09",x"c0",x"49"),
  1460 => (x"59",x"a6",x"f0",x"c0"),
  1461 => (x"48",x"66",x"ec",x"c0"),
  1462 => (x"c0",x"06",x"a8",x"c0"),
  1463 => (x"ec",x"c0",x"87",x"ee"),
  1464 => (x"a8",x"dd",x"48",x"66"),
  1465 => (x"87",x"e4",x"c0",x"03"),
  1466 => (x"49",x"bf",x"66",x"c4"),
  1467 => (x"81",x"66",x"ec",x"c0"),
  1468 => (x"c0",x"51",x"e0",x"c0"),
  1469 => (x"c1",x"49",x"66",x"ec"),
  1470 => (x"bf",x"66",x"c4",x"81"),
  1471 => (x"51",x"c1",x"c2",x"81"),
  1472 => (x"49",x"66",x"ec",x"c0"),
  1473 => (x"66",x"c4",x"81",x"c2"),
  1474 => (x"51",x"c0",x"81",x"bf"),
  1475 => (x"cc",x"c1",x"48",x"6e"),
  1476 => (x"49",x"6e",x"78",x"fd"),
  1477 => (x"66",x"d8",x"81",x"c8"),
  1478 => (x"c9",x"49",x"6e",x"51"),
  1479 => (x"51",x"66",x"d0",x"81"),
  1480 => (x"81",x"ca",x"49",x"6e"),
  1481 => (x"d8",x"51",x"66",x"dc"),
  1482 => (x"80",x"c1",x"48",x"66"),
  1483 => (x"48",x"58",x"a6",x"dc"),
  1484 => (x"78",x"c1",x"80",x"ec"),
  1485 => (x"ff",x"87",x"f2",x"c4"),
  1486 => (x"70",x"87",x"cb",x"dc"),
  1487 => (x"a6",x"f0",x"c0",x"49"),
  1488 => (x"c1",x"dc",x"ff",x"59"),
  1489 => (x"c0",x"49",x"70",x"87"),
  1490 => (x"dc",x"59",x"a6",x"e0"),
  1491 => (x"ec",x"c0",x"48",x"66"),
  1492 => (x"ca",x"c0",x"05",x"a8"),
  1493 => (x"48",x"a6",x"dc",x"87"),
  1494 => (x"78",x"66",x"ec",x"c0"),
  1495 => (x"ff",x"87",x"c4",x"c0"),
  1496 => (x"c8",x"87",x"cb",x"d8"),
  1497 => (x"91",x"cb",x"49",x"66"),
  1498 => (x"48",x"66",x"c4",x"c1"),
  1499 => (x"7e",x"70",x"80",x"71"),
  1500 => (x"82",x"c8",x"4a",x"6e"),
  1501 => (x"81",x"ca",x"49",x"6e"),
  1502 => (x"51",x"66",x"ec",x"c0"),
  1503 => (x"c1",x"49",x"66",x"dc"),
  1504 => (x"66",x"ec",x"c0",x"81"),
  1505 => (x"71",x"48",x"c1",x"89"),
  1506 => (x"c1",x"49",x"70",x"30"),
  1507 => (x"7a",x"97",x"71",x"89"),
  1508 => (x"bf",x"e0",x"f6",x"c2"),
  1509 => (x"66",x"ec",x"c0",x"49"),
  1510 => (x"4a",x"6a",x"97",x"29"),
  1511 => (x"c0",x"98",x"71",x"48"),
  1512 => (x"6e",x"58",x"a6",x"f4"),
  1513 => (x"a6",x"81",x"c4",x"49"),
  1514 => (x"c0",x"78",x"69",x"48"),
  1515 => (x"c0",x"48",x"66",x"e4"),
  1516 => (x"02",x"a8",x"66",x"e0"),
  1517 => (x"dc",x"87",x"c8",x"c0"),
  1518 => (x"78",x"c0",x"48",x"a6"),
  1519 => (x"dc",x"87",x"c5",x"c0"),
  1520 => (x"78",x"c1",x"48",x"a6"),
  1521 => (x"c0",x"1e",x"66",x"dc"),
  1522 => (x"66",x"cc",x"1e",x"e0"),
  1523 => (x"c6",x"d8",x"ff",x"49"),
  1524 => (x"70",x"86",x"c8",x"87"),
  1525 => (x"ac",x"b7",x"c0",x"4c"),
  1526 => (x"87",x"db",x"c1",x"06"),
  1527 => (x"74",x"48",x"66",x"c4"),
  1528 => (x"58",x"a6",x"c8",x"80"),
  1529 => (x"74",x"49",x"e0",x"c0"),
  1530 => (x"4b",x"66",x"c4",x"89"),
  1531 => (x"4a",x"ff",x"e3",x"c1"),
  1532 => (x"f3",x"e2",x"fe",x"71"),
  1533 => (x"48",x"66",x"c4",x"87"),
  1534 => (x"a6",x"c8",x"80",x"c2"),
  1535 => (x"66",x"e8",x"c0",x"58"),
  1536 => (x"c0",x"80",x"c1",x"48"),
  1537 => (x"c0",x"58",x"a6",x"ec"),
  1538 => (x"c1",x"49",x"66",x"f0"),
  1539 => (x"02",x"a9",x"70",x"81"),
  1540 => (x"c0",x"87",x"c5",x"c0"),
  1541 => (x"87",x"c2",x"c0",x"4d"),
  1542 => (x"1e",x"75",x"4d",x"c1"),
  1543 => (x"c0",x"49",x"a4",x"c2"),
  1544 => (x"88",x"71",x"48",x"e0"),
  1545 => (x"cc",x"1e",x"49",x"70"),
  1546 => (x"d6",x"ff",x"49",x"66"),
  1547 => (x"86",x"c8",x"87",x"e9"),
  1548 => (x"01",x"a8",x"b7",x"c0"),
  1549 => (x"c0",x"87",x"c6",x"ff"),
  1550 => (x"c0",x"02",x"66",x"e8"),
  1551 => (x"49",x"6e",x"87",x"d1"),
  1552 => (x"e8",x"c0",x"81",x"c9"),
  1553 => (x"48",x"6e",x"51",x"66"),
  1554 => (x"78",x"ce",x"cf",x"c1"),
  1555 => (x"6e",x"87",x"cc",x"c0"),
  1556 => (x"c2",x"81",x"c9",x"49"),
  1557 => (x"c1",x"48",x"6e",x"51"),
  1558 => (x"c4",x"78",x"c2",x"d0"),
  1559 => (x"78",x"c1",x"48",x"a6"),
  1560 => (x"ff",x"87",x"c6",x"c0"),
  1561 => (x"70",x"87",x"dc",x"d5"),
  1562 => (x"02",x"66",x"c4",x"4c"),
  1563 => (x"c8",x"87",x"f5",x"c0"),
  1564 => (x"66",x"cc",x"48",x"66"),
  1565 => (x"cb",x"c0",x"04",x"a8"),
  1566 => (x"48",x"66",x"c8",x"87"),
  1567 => (x"a6",x"cc",x"80",x"c1"),
  1568 => (x"87",x"e0",x"c0",x"58"),
  1569 => (x"c1",x"48",x"66",x"cc"),
  1570 => (x"58",x"a6",x"d0",x"88"),
  1571 => (x"c1",x"87",x"d5",x"c0"),
  1572 => (x"c0",x"05",x"ac",x"c6"),
  1573 => (x"66",x"d8",x"87",x"c8"),
  1574 => (x"dc",x"80",x"c1",x"48"),
  1575 => (x"d4",x"ff",x"58",x"a6"),
  1576 => (x"4c",x"70",x"87",x"e1"),
  1577 => (x"c1",x"48",x"66",x"d0"),
  1578 => (x"58",x"a6",x"d4",x"80"),
  1579 => (x"c0",x"02",x"9c",x"74"),
  1580 => (x"66",x"c8",x"87",x"cb"),
  1581 => (x"66",x"cc",x"c1",x"48"),
  1582 => (x"da",x"f3",x"04",x"a8"),
  1583 => (x"f9",x"d3",x"ff",x"87"),
  1584 => (x"48",x"66",x"c8",x"87"),
  1585 => (x"c0",x"03",x"a8",x"c7"),
  1586 => (x"f2",x"c2",x"87",x"e5"),
  1587 => (x"78",x"c0",x"48",x"f4"),
  1588 => (x"cb",x"49",x"66",x"c8"),
  1589 => (x"66",x"c4",x"c1",x"91"),
  1590 => (x"4a",x"a1",x"c4",x"81"),
  1591 => (x"52",x"c0",x"4a",x"6a"),
  1592 => (x"48",x"66",x"c8",x"79"),
  1593 => (x"a6",x"cc",x"80",x"c1"),
  1594 => (x"04",x"a8",x"c7",x"58"),
  1595 => (x"ff",x"87",x"db",x"ff"),
  1596 => (x"df",x"ff",x"8e",x"cc"),
  1597 => (x"6f",x"4c",x"87",x"f6"),
  1598 => (x"2a",x"20",x"64",x"61"),
  1599 => (x"3a",x"00",x"20",x"2e"),
  1600 => (x"49",x"44",x"00",x"20"),
  1601 => (x"77",x"53",x"20",x"50"),
  1602 => (x"68",x"63",x"74",x"69"),
  1603 => (x"1e",x"00",x"73",x"65"),
  1604 => (x"4b",x"71",x"1e",x"73"),
  1605 => (x"87",x"c6",x"02",x"9b"),
  1606 => (x"48",x"f0",x"f2",x"c2"),
  1607 => (x"1e",x"c7",x"78",x"c0"),
  1608 => (x"bf",x"f0",x"f2",x"c2"),
  1609 => (x"e7",x"c1",x"1e",x"49"),
  1610 => (x"f2",x"c2",x"1e",x"e4"),
  1611 => (x"ee",x"49",x"bf",x"d8"),
  1612 => (x"86",x"cc",x"87",x"c9"),
  1613 => (x"bf",x"d8",x"f2",x"c2"),
  1614 => (x"87",x"ea",x"e9",x"49"),
  1615 => (x"c8",x"02",x"9b",x"73"),
  1616 => (x"e4",x"e7",x"c1",x"87"),
  1617 => (x"e6",x"ed",x"c0",x"49"),
  1618 => (x"e3",x"de",x"ff",x"87"),
  1619 => (x"cd",x"c7",x"1e",x"87"),
  1620 => (x"fe",x"49",x"c1",x"87"),
  1621 => (x"e5",x"fe",x"87",x"f9"),
  1622 => (x"98",x"70",x"87",x"dc"),
  1623 => (x"fe",x"87",x"cd",x"02"),
  1624 => (x"70",x"87",x"f5",x"ec"),
  1625 => (x"87",x"c4",x"02",x"98"),
  1626 => (x"87",x"c2",x"4a",x"c1"),
  1627 => (x"9a",x"72",x"4a",x"c0"),
  1628 => (x"c0",x"87",x"ce",x"05"),
  1629 => (x"e2",x"e6",x"c1",x"1e"),
  1630 => (x"d0",x"f9",x"c0",x"49"),
  1631 => (x"fe",x"86",x"c4",x"87"),
  1632 => (x"f3",x"fb",x"c0",x"87"),
  1633 => (x"c1",x"1e",x"c0",x"87"),
  1634 => (x"c0",x"49",x"ed",x"e6"),
  1635 => (x"c0",x"87",x"fe",x"f8"),
  1636 => (x"f9",x"fd",x"c0",x"1e"),
  1637 => (x"c0",x"49",x"70",x"87"),
  1638 => (x"c2",x"87",x"f2",x"f8"),
  1639 => (x"8e",x"f8",x"87",x"ff"),
  1640 => (x"44",x"53",x"4f",x"26"),
  1641 => (x"69",x"61",x"66",x"20"),
  1642 => (x"2e",x"64",x"65",x"6c"),
  1643 => (x"6f",x"6f",x"42",x"00"),
  1644 => (x"67",x"6e",x"69",x"74"),
  1645 => (x"00",x"2e",x"2e",x"2e"),
  1646 => (x"f0",x"f2",x"c2",x"1e"),
  1647 => (x"c2",x"78",x"c0",x"48"),
  1648 => (x"c0",x"48",x"d8",x"f2"),
  1649 => (x"87",x"c5",x"fe",x"78"),
  1650 => (x"87",x"e1",x"fd",x"c0"),
  1651 => (x"4f",x"26",x"48",x"c0"),
  1652 => (x"00",x"01",x"00",x"00"),
  1653 => (x"20",x"80",x"00",x"00"),
  1654 => (x"74",x"69",x"78",x"45"),
  1655 => (x"42",x"20",x"80",x"00"),
  1656 => (x"00",x"6b",x"63",x"61"),
  1657 => (x"00",x"00",x"13",x"7e"),
  1658 => (x"00",x"00",x"2c",x"c4"),
  1659 => (x"7e",x"00",x"00",x"00"),
  1660 => (x"e2",x"00",x"00",x"13"),
  1661 => (x"00",x"00",x"00",x"2c"),
  1662 => (x"13",x"7e",x"00",x"00"),
  1663 => (x"2d",x"00",x"00",x"00"),
  1664 => (x"00",x"00",x"00",x"00"),
  1665 => (x"00",x"13",x"7e",x"00"),
  1666 => (x"00",x"2d",x"1e",x"00"),
  1667 => (x"00",x"00",x"00",x"00"),
  1668 => (x"00",x"00",x"13",x"7e"),
  1669 => (x"00",x"00",x"2d",x"3c"),
  1670 => (x"7e",x"00",x"00",x"00"),
  1671 => (x"5a",x"00",x"00",x"13"),
  1672 => (x"00",x"00",x"00",x"2d"),
  1673 => (x"13",x"7e",x"00",x"00"),
  1674 => (x"2d",x"78",x"00",x"00"),
  1675 => (x"00",x"00",x"00",x"00"),
  1676 => (x"00",x"13",x"7e",x"00"),
  1677 => (x"00",x"00",x"00",x"00"),
  1678 => (x"00",x"00",x"00",x"00"),
  1679 => (x"00",x"00",x"14",x"13"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"1e",x"00",x"00",x"00"),
  1682 => (x"c0",x"48",x"f0",x"fe"),
  1683 => (x"79",x"09",x"cd",x"78"),
  1684 => (x"1e",x"4f",x"26",x"09"),
  1685 => (x"bf",x"f0",x"fe",x"1e"),
  1686 => (x"26",x"26",x"48",x"7e"),
  1687 => (x"f0",x"fe",x"1e",x"4f"),
  1688 => (x"26",x"78",x"c1",x"48"),
  1689 => (x"f0",x"fe",x"1e",x"4f"),
  1690 => (x"26",x"78",x"c0",x"48"),
  1691 => (x"4a",x"71",x"1e",x"4f"),
  1692 => (x"26",x"52",x"52",x"c0"),
  1693 => (x"5b",x"5e",x"0e",x"4f"),
  1694 => (x"f4",x"0e",x"5d",x"5c"),
  1695 => (x"97",x"4d",x"71",x"86"),
  1696 => (x"a5",x"c1",x"7e",x"6d"),
  1697 => (x"48",x"6c",x"97",x"4c"),
  1698 => (x"6e",x"58",x"a6",x"c8"),
  1699 => (x"a8",x"66",x"c4",x"48"),
  1700 => (x"ff",x"87",x"c5",x"05"),
  1701 => (x"87",x"e6",x"c0",x"48"),
  1702 => (x"c2",x"87",x"ca",x"ff"),
  1703 => (x"6c",x"97",x"49",x"a5"),
  1704 => (x"4b",x"a3",x"71",x"4b"),
  1705 => (x"97",x"4b",x"6b",x"97"),
  1706 => (x"48",x"6e",x"7e",x"6c"),
  1707 => (x"a6",x"c8",x"80",x"c1"),
  1708 => (x"cc",x"98",x"c7",x"58"),
  1709 => (x"97",x"70",x"58",x"a6"),
  1710 => (x"87",x"e1",x"fe",x"7c"),
  1711 => (x"8e",x"f4",x"48",x"73"),
  1712 => (x"4c",x"26",x"4d",x"26"),
  1713 => (x"4f",x"26",x"4b",x"26"),
  1714 => (x"5c",x"5b",x"5e",x"0e"),
  1715 => (x"71",x"86",x"f4",x"0e"),
  1716 => (x"4a",x"66",x"d8",x"4c"),
  1717 => (x"c2",x"9a",x"ff",x"c3"),
  1718 => (x"6c",x"97",x"4b",x"a4"),
  1719 => (x"49",x"a1",x"73",x"49"),
  1720 => (x"6c",x"97",x"51",x"72"),
  1721 => (x"c1",x"48",x"6e",x"7e"),
  1722 => (x"58",x"a6",x"c8",x"80"),
  1723 => (x"a6",x"cc",x"98",x"c7"),
  1724 => (x"f4",x"54",x"70",x"58"),
  1725 => (x"87",x"ca",x"ff",x"8e"),
  1726 => (x"e8",x"fd",x"1e",x"1e"),
  1727 => (x"4a",x"bf",x"e0",x"87"),
  1728 => (x"c0",x"e0",x"c0",x"49"),
  1729 => (x"87",x"cb",x"02",x"99"),
  1730 => (x"f6",x"c2",x"1e",x"72"),
  1731 => (x"f7",x"fe",x"49",x"d6"),
  1732 => (x"fc",x"86",x"c4",x"87"),
  1733 => (x"7e",x"70",x"87",x"fd"),
  1734 => (x"26",x"87",x"c2",x"fd"),
  1735 => (x"c2",x"1e",x"4f",x"26"),
  1736 => (x"fd",x"49",x"d6",x"f6"),
  1737 => (x"eb",x"c1",x"87",x"c7"),
  1738 => (x"da",x"fc",x"49",x"f8"),
  1739 => (x"87",x"c7",x"c4",x"87"),
  1740 => (x"ff",x"1e",x"4f",x"26"),
  1741 => (x"e1",x"c8",x"48",x"d0"),
  1742 => (x"48",x"d4",x"ff",x"78"),
  1743 => (x"66",x"c4",x"78",x"c5"),
  1744 => (x"c3",x"87",x"c3",x"02"),
  1745 => (x"66",x"c8",x"78",x"e0"),
  1746 => (x"ff",x"87",x"c6",x"02"),
  1747 => (x"f0",x"c3",x"48",x"d4"),
  1748 => (x"48",x"d4",x"ff",x"78"),
  1749 => (x"d0",x"ff",x"78",x"71"),
  1750 => (x"78",x"e1",x"c8",x"48"),
  1751 => (x"26",x"78",x"e0",x"c0"),
  1752 => (x"5b",x"5e",x"0e",x"4f"),
  1753 => (x"4c",x"71",x"0e",x"5c"),
  1754 => (x"49",x"d6",x"f6",x"c2"),
  1755 => (x"70",x"87",x"c6",x"fc"),
  1756 => (x"aa",x"b7",x"c0",x"4a"),
  1757 => (x"87",x"e2",x"c2",x"04"),
  1758 => (x"05",x"aa",x"f0",x"c3"),
  1759 => (x"f0",x"c1",x"87",x"c9"),
  1760 => (x"78",x"c1",x"48",x"e6"),
  1761 => (x"c3",x"87",x"c3",x"c2"),
  1762 => (x"c9",x"05",x"aa",x"e0"),
  1763 => (x"ea",x"f0",x"c1",x"87"),
  1764 => (x"c1",x"78",x"c1",x"48"),
  1765 => (x"f0",x"c1",x"87",x"f4"),
  1766 => (x"c6",x"02",x"bf",x"ea"),
  1767 => (x"a2",x"c0",x"c2",x"87"),
  1768 => (x"72",x"87",x"c2",x"4b"),
  1769 => (x"05",x"9c",x"74",x"4b"),
  1770 => (x"f0",x"c1",x"87",x"d1"),
  1771 => (x"c1",x"1e",x"bf",x"e6"),
  1772 => (x"1e",x"bf",x"ea",x"f0"),
  1773 => (x"f9",x"fd",x"49",x"72"),
  1774 => (x"c1",x"86",x"c8",x"87"),
  1775 => (x"02",x"bf",x"e6",x"f0"),
  1776 => (x"73",x"87",x"e0",x"c0"),
  1777 => (x"29",x"b7",x"c4",x"49"),
  1778 => (x"c6",x"f2",x"c1",x"91"),
  1779 => (x"cf",x"4a",x"73",x"81"),
  1780 => (x"c1",x"92",x"c2",x"9a"),
  1781 => (x"70",x"30",x"72",x"48"),
  1782 => (x"72",x"ba",x"ff",x"4a"),
  1783 => (x"70",x"98",x"69",x"48"),
  1784 => (x"73",x"87",x"db",x"79"),
  1785 => (x"29",x"b7",x"c4",x"49"),
  1786 => (x"c6",x"f2",x"c1",x"91"),
  1787 => (x"cf",x"4a",x"73",x"81"),
  1788 => (x"c3",x"92",x"c2",x"9a"),
  1789 => (x"70",x"30",x"72",x"48"),
  1790 => (x"b0",x"69",x"48",x"4a"),
  1791 => (x"f0",x"c1",x"79",x"70"),
  1792 => (x"78",x"c0",x"48",x"ea"),
  1793 => (x"48",x"e6",x"f0",x"c1"),
  1794 => (x"f6",x"c2",x"78",x"c0"),
  1795 => (x"e4",x"f9",x"49",x"d6"),
  1796 => (x"c0",x"4a",x"70",x"87"),
  1797 => (x"fd",x"03",x"aa",x"b7"),
  1798 => (x"48",x"c0",x"87",x"de"),
  1799 => (x"4d",x"26",x"87",x"c2"),
  1800 => (x"4b",x"26",x"4c",x"26"),
  1801 => (x"00",x"00",x"4f",x"26"),
  1802 => (x"00",x"00",x"00",x"00"),
  1803 => (x"71",x"1e",x"00",x"00"),
  1804 => (x"ec",x"fc",x"49",x"4a"),
  1805 => (x"1e",x"4f",x"26",x"87"),
  1806 => (x"49",x"72",x"4a",x"c0"),
  1807 => (x"f2",x"c1",x"91",x"c4"),
  1808 => (x"79",x"c0",x"81",x"c6"),
  1809 => (x"b7",x"d0",x"82",x"c1"),
  1810 => (x"87",x"ee",x"04",x"aa"),
  1811 => (x"5e",x"0e",x"4f",x"26"),
  1812 => (x"0e",x"5d",x"5c",x"5b"),
  1813 => (x"cc",x"f8",x"4d",x"71"),
  1814 => (x"c4",x"4a",x"75",x"87"),
  1815 => (x"c1",x"92",x"2a",x"b7"),
  1816 => (x"75",x"82",x"c6",x"f2"),
  1817 => (x"c2",x"9c",x"cf",x"4c"),
  1818 => (x"4b",x"49",x"6a",x"94"),
  1819 => (x"9b",x"c3",x"2b",x"74"),
  1820 => (x"30",x"74",x"48",x"c2"),
  1821 => (x"bc",x"ff",x"4c",x"70"),
  1822 => (x"98",x"71",x"48",x"74"),
  1823 => (x"dc",x"f7",x"7a",x"70"),
  1824 => (x"fe",x"48",x"73",x"87"),
  1825 => (x"00",x"00",x"87",x"d8"),
  1826 => (x"00",x"00",x"00",x"00"),
  1827 => (x"00",x"00",x"00",x"00"),
  1828 => (x"00",x"00",x"00",x"00"),
  1829 => (x"00",x"00",x"00",x"00"),
  1830 => (x"00",x"00",x"00",x"00"),
  1831 => (x"00",x"00",x"00",x"00"),
  1832 => (x"00",x"00",x"00",x"00"),
  1833 => (x"00",x"00",x"00",x"00"),
  1834 => (x"00",x"00",x"00",x"00"),
  1835 => (x"00",x"00",x"00",x"00"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"00",x"00",x"00",x"00"),
  1838 => (x"00",x"00",x"00",x"00"),
  1839 => (x"00",x"00",x"00",x"00"),
  1840 => (x"00",x"00",x"00",x"00"),
  1841 => (x"ff",x"1e",x"00",x"00"),
  1842 => (x"e1",x"c8",x"48",x"d0"),
  1843 => (x"ff",x"48",x"71",x"78"),
  1844 => (x"c4",x"78",x"08",x"d4"),
  1845 => (x"d4",x"ff",x"48",x"66"),
  1846 => (x"4f",x"26",x"78",x"08"),
  1847 => (x"c4",x"4a",x"71",x"1e"),
  1848 => (x"72",x"1e",x"49",x"66"),
  1849 => (x"87",x"de",x"ff",x"49"),
  1850 => (x"c0",x"48",x"d0",x"ff"),
  1851 => (x"26",x"26",x"78",x"e0"),
  1852 => (x"1e",x"73",x"1e",x"4f"),
  1853 => (x"66",x"c8",x"4b",x"71"),
  1854 => (x"4a",x"73",x"1e",x"49"),
  1855 => (x"49",x"a2",x"e0",x"c1"),
  1856 => (x"26",x"87",x"d9",x"ff"),
  1857 => (x"4d",x"26",x"87",x"c4"),
  1858 => (x"4b",x"26",x"4c",x"26"),
  1859 => (x"ff",x"1e",x"4f",x"26"),
  1860 => (x"ff",x"c3",x"4a",x"d4"),
  1861 => (x"48",x"d0",x"ff",x"7a"),
  1862 => (x"de",x"78",x"e1",x"c0"),
  1863 => (x"e0",x"f6",x"c2",x"7a"),
  1864 => (x"48",x"49",x"7a",x"bf"),
  1865 => (x"7a",x"70",x"28",x"c8"),
  1866 => (x"28",x"d0",x"48",x"71"),
  1867 => (x"48",x"71",x"7a",x"70"),
  1868 => (x"7a",x"70",x"28",x"d8"),
  1869 => (x"c0",x"48",x"d0",x"ff"),
  1870 => (x"4f",x"26",x"78",x"e0"),
  1871 => (x"5c",x"5b",x"5e",x"0e"),
  1872 => (x"4c",x"71",x"0e",x"5d"),
  1873 => (x"bf",x"e0",x"f6",x"c2"),
  1874 => (x"2b",x"74",x"4b",x"4d"),
  1875 => (x"c1",x"9b",x"66",x"d0"),
  1876 => (x"ab",x"66",x"d4",x"83"),
  1877 => (x"c0",x"87",x"c2",x"04"),
  1878 => (x"d0",x"4a",x"74",x"4b"),
  1879 => (x"31",x"72",x"49",x"66"),
  1880 => (x"99",x"75",x"b9",x"ff"),
  1881 => (x"30",x"72",x"48",x"73"),
  1882 => (x"71",x"48",x"4a",x"70"),
  1883 => (x"e4",x"f6",x"c2",x"b0"),
  1884 => (x"87",x"da",x"fe",x"58"),
  1885 => (x"4c",x"26",x"4d",x"26"),
  1886 => (x"4f",x"26",x"4b",x"26"),
  1887 => (x"5c",x"5b",x"5e",x"0e"),
  1888 => (x"71",x"1e",x"0e",x"5d"),
  1889 => (x"e4",x"f6",x"c2",x"4c"),
  1890 => (x"c0",x"4a",x"c0",x"4b"),
  1891 => (x"cc",x"fe",x"49",x"f4"),
  1892 => (x"1e",x"74",x"87",x"e6"),
  1893 => (x"49",x"e4",x"f6",x"c2"),
  1894 => (x"87",x"e9",x"e7",x"fe"),
  1895 => (x"49",x"70",x"86",x"c4"),
  1896 => (x"ea",x"c0",x"02",x"99"),
  1897 => (x"a6",x"1e",x"c4",x"87"),
  1898 => (x"f6",x"c2",x"1e",x"4d"),
  1899 => (x"ef",x"fe",x"49",x"e4"),
  1900 => (x"86",x"c8",x"87",x"c0"),
  1901 => (x"d6",x"02",x"98",x"70"),
  1902 => (x"c1",x"4a",x"75",x"87"),
  1903 => (x"c4",x"49",x"c5",x"f8"),
  1904 => (x"e5",x"ca",x"fe",x"4b"),
  1905 => (x"02",x"98",x"70",x"87"),
  1906 => (x"48",x"c0",x"87",x"ca"),
  1907 => (x"c0",x"87",x"ed",x"c0"),
  1908 => (x"87",x"e8",x"c0",x"48"),
  1909 => (x"c1",x"87",x"f3",x"c0"),
  1910 => (x"98",x"70",x"87",x"c4"),
  1911 => (x"c0",x"87",x"c8",x"02"),
  1912 => (x"98",x"70",x"87",x"fc"),
  1913 => (x"c2",x"87",x"f8",x"05"),
  1914 => (x"02",x"bf",x"c4",x"f7"),
  1915 => (x"f6",x"c2",x"87",x"cc"),
  1916 => (x"f7",x"c2",x"48",x"e0"),
  1917 => (x"fc",x"78",x"bf",x"c4"),
  1918 => (x"48",x"c1",x"87",x"d4"),
  1919 => (x"26",x"4d",x"26",x"26"),
  1920 => (x"26",x"4b",x"26",x"4c"),
  1921 => (x"52",x"41",x"5b",x"4f"),
  1922 => (x"c0",x"1e",x"00",x"43"),
  1923 => (x"e4",x"f6",x"c2",x"1e"),
  1924 => (x"f2",x"eb",x"fe",x"49"),
  1925 => (x"fc",x"f6",x"c2",x"87"),
  1926 => (x"26",x"78",x"c0",x"48"),
  1927 => (x"5e",x"0e",x"4f",x"26"),
  1928 => (x"0e",x"5d",x"5c",x"5b"),
  1929 => (x"7e",x"c0",x"86",x"f4"),
  1930 => (x"bf",x"fc",x"f6",x"c2"),
  1931 => (x"a8",x"b7",x"c3",x"48"),
  1932 => (x"c2",x"87",x"d1",x"03"),
  1933 => (x"48",x"bf",x"fc",x"f6"),
  1934 => (x"f7",x"c2",x"80",x"c1"),
  1935 => (x"fb",x"c0",x"58",x"c0"),
  1936 => (x"87",x"d9",x"c6",x"48"),
  1937 => (x"49",x"e4",x"f6",x"c2"),
  1938 => (x"87",x"fa",x"f0",x"fe"),
  1939 => (x"b7",x"c0",x"4c",x"70"),
  1940 => (x"87",x"c4",x"03",x"ac"),
  1941 => (x"87",x"c5",x"c6",x"48"),
  1942 => (x"bf",x"fc",x"f6",x"c2"),
  1943 => (x"02",x"8a",x"c3",x"4a"),
  1944 => (x"8a",x"c1",x"87",x"d8"),
  1945 => (x"87",x"c7",x"c5",x"02"),
  1946 => (x"f2",x"c2",x"02",x"8a"),
  1947 => (x"c1",x"02",x"8a",x"87"),
  1948 => (x"02",x"8a",x"87",x"cf"),
  1949 => (x"c5",x"87",x"de",x"c3"),
  1950 => (x"4d",x"c0",x"87",x"d9"),
  1951 => (x"75",x"5c",x"a6",x"c8"),
  1952 => (x"c1",x"92",x"c4",x"4a"),
  1953 => (x"c2",x"82",x"fb",x"ff"),
  1954 => (x"75",x"4c",x"f8",x"f6"),
  1955 => (x"4b",x"6c",x"97",x"84"),
  1956 => (x"a3",x"c1",x"4b",x"49"),
  1957 => (x"81",x"6a",x"7c",x"97"),
  1958 => (x"a6",x"cc",x"48",x"11"),
  1959 => (x"48",x"66",x"c4",x"58"),
  1960 => (x"02",x"a8",x"66",x"c8"),
  1961 => (x"97",x"c0",x"87",x"c3"),
  1962 => (x"05",x"66",x"c8",x"7c"),
  1963 => (x"f6",x"c2",x"87",x"c7"),
  1964 => (x"a5",x"c4",x"48",x"fc"),
  1965 => (x"c4",x"85",x"c1",x"78"),
  1966 => (x"ff",x"04",x"ad",x"b7"),
  1967 => (x"d2",x"c4",x"87",x"c1"),
  1968 => (x"c8",x"f7",x"c2",x"87"),
  1969 => (x"b7",x"c8",x"48",x"bf"),
  1970 => (x"87",x"cb",x"01",x"a8"),
  1971 => (x"c6",x"02",x"ac",x"ca"),
  1972 => (x"05",x"ac",x"cd",x"87"),
  1973 => (x"c2",x"87",x"f3",x"c0"),
  1974 => (x"4b",x"bf",x"c8",x"f7"),
  1975 => (x"03",x"ab",x"b7",x"c8"),
  1976 => (x"f7",x"c2",x"87",x"d2"),
  1977 => (x"81",x"73",x"49",x"cc"),
  1978 => (x"c1",x"51",x"e0",x"c0"),
  1979 => (x"ab",x"b7",x"c8",x"83"),
  1980 => (x"87",x"ee",x"ff",x"04"),
  1981 => (x"48",x"d4",x"f7",x"c2"),
  1982 => (x"c1",x"50",x"d2",x"c1"),
  1983 => (x"cd",x"c1",x"50",x"cf"),
  1984 => (x"e4",x"50",x"c0",x"50"),
  1985 => (x"c3",x"78",x"c3",x"80"),
  1986 => (x"f7",x"c2",x"87",x"c9"),
  1987 => (x"48",x"49",x"bf",x"c8"),
  1988 => (x"f7",x"c2",x"80",x"c1"),
  1989 => (x"c4",x"48",x"58",x"cc"),
  1990 => (x"51",x"74",x"81",x"a0"),
  1991 => (x"c0",x"87",x"f4",x"c2"),
  1992 => (x"04",x"ac",x"b7",x"f0"),
  1993 => (x"f9",x"c0",x"87",x"da"),
  1994 => (x"d3",x"01",x"ac",x"b7"),
  1995 => (x"c0",x"f7",x"c2",x"87"),
  1996 => (x"91",x"ca",x"49",x"bf"),
  1997 => (x"f0",x"c0",x"4a",x"74"),
  1998 => (x"c0",x"f7",x"c2",x"8a"),
  1999 => (x"78",x"a1",x"72",x"48"),
  2000 => (x"c0",x"02",x"ac",x"ca"),
  2001 => (x"ac",x"cd",x"87",x"c6"),
  2002 => (x"87",x"c7",x"c2",x"05"),
  2003 => (x"48",x"fc",x"f6",x"c2"),
  2004 => (x"fe",x"c1",x"78",x"c3"),
  2005 => (x"b7",x"f0",x"c0",x"87"),
  2006 => (x"87",x"db",x"04",x"ac"),
  2007 => (x"ac",x"b7",x"f9",x"c0"),
  2008 => (x"87",x"d3",x"c0",x"01"),
  2009 => (x"bf",x"c4",x"f7",x"c2"),
  2010 => (x"74",x"91",x"d0",x"49"),
  2011 => (x"8a",x"f0",x"c0",x"4a"),
  2012 => (x"48",x"c4",x"f7",x"c2"),
  2013 => (x"c1",x"78",x"a1",x"72"),
  2014 => (x"04",x"ac",x"b7",x"c1"),
  2015 => (x"c1",x"87",x"db",x"c0"),
  2016 => (x"01",x"ac",x"b7",x"c6"),
  2017 => (x"c2",x"87",x"d3",x"c0"),
  2018 => (x"49",x"bf",x"c4",x"f7"),
  2019 => (x"4a",x"74",x"91",x"d0"),
  2020 => (x"c2",x"8a",x"f7",x"c0"),
  2021 => (x"72",x"48",x"c4",x"f7"),
  2022 => (x"ac",x"ca",x"78",x"a1"),
  2023 => (x"87",x"c6",x"c0",x"02"),
  2024 => (x"c0",x"05",x"ac",x"cd"),
  2025 => (x"f6",x"c2",x"87",x"ed"),
  2026 => (x"78",x"c3",x"48",x"fc"),
  2027 => (x"c0",x"87",x"e4",x"c0"),
  2028 => (x"c0",x"05",x"ac",x"e2"),
  2029 => (x"fb",x"c0",x"87",x"c6"),
  2030 => (x"87",x"d7",x"c0",x"7e"),
  2031 => (x"c0",x"02",x"ac",x"ca"),
  2032 => (x"ac",x"cd",x"87",x"c6"),
  2033 => (x"87",x"c9",x"c0",x"05"),
  2034 => (x"48",x"fc",x"f6",x"c2"),
  2035 => (x"c2",x"c0",x"78",x"c3"),
  2036 => (x"6e",x"7e",x"74",x"87"),
  2037 => (x"87",x"d0",x"f9",x"02"),
  2038 => (x"ff",x"c3",x"48",x"6e"),
  2039 => (x"f8",x"8e",x"f4",x"99"),
  2040 => (x"4f",x"43",x"87",x"db"),
  2041 => (x"00",x"3d",x"46",x"4e"),
  2042 => (x"00",x"44",x"4f",x"4d"),
  2043 => (x"45",x"4d",x"41",x"4e"),
  2044 => (x"46",x"45",x"44",x"00"),
  2045 => (x"54",x"4c",x"55",x"41"),
  2046 => (x"e2",x"00",x"30",x"3d"),
  2047 => (x"e8",x"00",x"00",x"1f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

