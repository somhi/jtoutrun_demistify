
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"45",x"4d",x"41",x"4e"),
     1 => (x"46",x"45",x"44",x"00"),
     2 => (x"54",x"4c",x"55",x"41"),
     3 => (x"f6",x"00",x"30",x"3d"),
     4 => (x"fc",x"00",x"00",x"1f"),
     5 => (x"00",x"00",x"00",x"1f"),
     6 => (x"05",x"00",x"00",x"20"),
     7 => (x"1e",x"00",x"00",x"20"),
     8 => (x"c8",x"48",x"d0",x"ff"),
     9 => (x"48",x"71",x"78",x"c9"),
    10 => (x"78",x"08",x"d4",x"ff"),
    11 => (x"71",x"1e",x"4f",x"26"),
    12 => (x"87",x"eb",x"49",x"4a"),
    13 => (x"c8",x"48",x"d0",x"ff"),
    14 => (x"1e",x"4f",x"26",x"78"),
    15 => (x"4b",x"71",x"1e",x"73"),
    16 => (x"bf",x"f8",x"f7",x"c2"),
    17 => (x"c2",x"87",x"c3",x"02"),
    18 => (x"d0",x"ff",x"87",x"eb"),
    19 => (x"78",x"c9",x"c8",x"48"),
    20 => (x"e0",x"c0",x"49",x"73"),
    21 => (x"48",x"d4",x"ff",x"b1"),
    22 => (x"f7",x"c2",x"78",x"71"),
    23 => (x"78",x"c0",x"48",x"ec"),
    24 => (x"c5",x"02",x"66",x"c8"),
    25 => (x"49",x"ff",x"c3",x"87"),
    26 => (x"49",x"c0",x"87",x"c2"),
    27 => (x"59",x"f4",x"f7",x"c2"),
    28 => (x"c6",x"02",x"66",x"cc"),
    29 => (x"d5",x"d5",x"c5",x"87"),
    30 => (x"cf",x"87",x"c4",x"4a"),
    31 => (x"c2",x"4a",x"ff",x"ff"),
    32 => (x"c2",x"5a",x"f8",x"f7"),
    33 => (x"c1",x"48",x"f8",x"f7"),
    34 => (x"26",x"87",x"c4",x"78"),
    35 => (x"26",x"4c",x"26",x"4d"),
    36 => (x"0e",x"4f",x"26",x"4b"),
    37 => (x"5d",x"5c",x"5b",x"5e"),
    38 => (x"c2",x"4a",x"71",x"0e"),
    39 => (x"4c",x"bf",x"f4",x"f7"),
    40 => (x"cb",x"02",x"9a",x"72"),
    41 => (x"91",x"c8",x"49",x"87"),
    42 => (x"4b",x"f1",x"c0",x"c2"),
    43 => (x"87",x"c4",x"83",x"71"),
    44 => (x"4b",x"f1",x"c4",x"c2"),
    45 => (x"49",x"13",x"4d",x"c0"),
    46 => (x"f7",x"c2",x"99",x"74"),
    47 => (x"ff",x"b9",x"bf",x"f0"),
    48 => (x"78",x"71",x"48",x"d4"),
    49 => (x"85",x"2c",x"b7",x"c1"),
    50 => (x"04",x"ad",x"b7",x"c8"),
    51 => (x"f7",x"c2",x"87",x"e8"),
    52 => (x"c8",x"48",x"bf",x"ec"),
    53 => (x"f0",x"f7",x"c2",x"80"),
    54 => (x"87",x"ef",x"fe",x"58"),
    55 => (x"71",x"1e",x"73",x"1e"),
    56 => (x"9a",x"4a",x"13",x"4b"),
    57 => (x"72",x"87",x"cb",x"02"),
    58 => (x"87",x"e7",x"fe",x"49"),
    59 => (x"05",x"9a",x"4a",x"13"),
    60 => (x"da",x"fe",x"87",x"f5"),
    61 => (x"f7",x"c2",x"1e",x"87"),
    62 => (x"c2",x"49",x"bf",x"ec"),
    63 => (x"c1",x"48",x"ec",x"f7"),
    64 => (x"c0",x"c4",x"78",x"a1"),
    65 => (x"db",x"03",x"a9",x"b7"),
    66 => (x"48",x"d4",x"ff",x"87"),
    67 => (x"bf",x"f0",x"f7",x"c2"),
    68 => (x"ec",x"f7",x"c2",x"78"),
    69 => (x"f7",x"c2",x"49",x"bf"),
    70 => (x"a1",x"c1",x"48",x"ec"),
    71 => (x"b7",x"c0",x"c4",x"78"),
    72 => (x"87",x"e5",x"04",x"a9"),
    73 => (x"c8",x"48",x"d0",x"ff"),
    74 => (x"f8",x"f7",x"c2",x"78"),
    75 => (x"26",x"78",x"c0",x"48"),
    76 => (x"00",x"00",x"00",x"4f"),
    77 => (x"00",x"00",x"00",x"00"),
    78 => (x"00",x"00",x"00",x"00"),
    79 => (x"00",x"00",x"5f",x"5f"),
    80 => (x"03",x"03",x"00",x"00"),
    81 => (x"00",x"03",x"03",x"00"),
    82 => (x"7f",x"7f",x"14",x"00"),
    83 => (x"14",x"7f",x"7f",x"14"),
    84 => (x"2e",x"24",x"00",x"00"),
    85 => (x"12",x"3a",x"6b",x"6b"),
    86 => (x"36",x"6a",x"4c",x"00"),
    87 => (x"32",x"56",x"6c",x"18"),
    88 => (x"4f",x"7e",x"30",x"00"),
    89 => (x"68",x"3a",x"77",x"59"),
    90 => (x"04",x"00",x"00",x"40"),
    91 => (x"00",x"00",x"03",x"07"),
    92 => (x"1c",x"00",x"00",x"00"),
    93 => (x"00",x"41",x"63",x"3e"),
    94 => (x"41",x"00",x"00",x"00"),
    95 => (x"00",x"1c",x"3e",x"63"),
    96 => (x"3e",x"2a",x"08",x"00"),
    97 => (x"2a",x"3e",x"1c",x"1c"),
    98 => (x"08",x"08",x"00",x"08"),
    99 => (x"08",x"08",x"3e",x"3e"),
   100 => (x"80",x"00",x"00",x"00"),
   101 => (x"00",x"00",x"60",x"e0"),
   102 => (x"08",x"08",x"00",x"00"),
   103 => (x"08",x"08",x"08",x"08"),
   104 => (x"00",x"00",x"00",x"00"),
   105 => (x"00",x"00",x"60",x"60"),
   106 => (x"30",x"60",x"40",x"00"),
   107 => (x"03",x"06",x"0c",x"18"),
   108 => (x"7f",x"3e",x"00",x"01"),
   109 => (x"3e",x"7f",x"4d",x"59"),
   110 => (x"06",x"04",x"00",x"00"),
   111 => (x"00",x"00",x"7f",x"7f"),
   112 => (x"63",x"42",x"00",x"00"),
   113 => (x"46",x"4f",x"59",x"71"),
   114 => (x"63",x"22",x"00",x"00"),
   115 => (x"36",x"7f",x"49",x"49"),
   116 => (x"16",x"1c",x"18",x"00"),
   117 => (x"10",x"7f",x"7f",x"13"),
   118 => (x"67",x"27",x"00",x"00"),
   119 => (x"39",x"7d",x"45",x"45"),
   120 => (x"7e",x"3c",x"00",x"00"),
   121 => (x"30",x"79",x"49",x"4b"),
   122 => (x"01",x"01",x"00",x"00"),
   123 => (x"07",x"0f",x"79",x"71"),
   124 => (x"7f",x"36",x"00",x"00"),
   125 => (x"36",x"7f",x"49",x"49"),
   126 => (x"4f",x"06",x"00",x"00"),
   127 => (x"1e",x"3f",x"69",x"49"),
   128 => (x"00",x"00",x"00",x"00"),
   129 => (x"00",x"00",x"66",x"66"),
   130 => (x"80",x"00",x"00",x"00"),
   131 => (x"00",x"00",x"66",x"e6"),
   132 => (x"08",x"08",x"00",x"00"),
   133 => (x"22",x"22",x"14",x"14"),
   134 => (x"14",x"14",x"00",x"00"),
   135 => (x"14",x"14",x"14",x"14"),
   136 => (x"22",x"22",x"00",x"00"),
   137 => (x"08",x"08",x"14",x"14"),
   138 => (x"03",x"02",x"00",x"00"),
   139 => (x"06",x"0f",x"59",x"51"),
   140 => (x"41",x"7f",x"3e",x"00"),
   141 => (x"1e",x"1f",x"55",x"5d"),
   142 => (x"7f",x"7e",x"00",x"00"),
   143 => (x"7e",x"7f",x"09",x"09"),
   144 => (x"7f",x"7f",x"00",x"00"),
   145 => (x"36",x"7f",x"49",x"49"),
   146 => (x"3e",x"1c",x"00",x"00"),
   147 => (x"41",x"41",x"41",x"63"),
   148 => (x"7f",x"7f",x"00",x"00"),
   149 => (x"1c",x"3e",x"63",x"41"),
   150 => (x"7f",x"7f",x"00",x"00"),
   151 => (x"41",x"41",x"49",x"49"),
   152 => (x"7f",x"7f",x"00",x"00"),
   153 => (x"01",x"01",x"09",x"09"),
   154 => (x"7f",x"3e",x"00",x"00"),
   155 => (x"7a",x"7b",x"49",x"41"),
   156 => (x"7f",x"7f",x"00",x"00"),
   157 => (x"7f",x"7f",x"08",x"08"),
   158 => (x"41",x"00",x"00",x"00"),
   159 => (x"00",x"41",x"7f",x"7f"),
   160 => (x"60",x"20",x"00",x"00"),
   161 => (x"3f",x"7f",x"40",x"40"),
   162 => (x"08",x"7f",x"7f",x"00"),
   163 => (x"41",x"63",x"36",x"1c"),
   164 => (x"7f",x"7f",x"00",x"00"),
   165 => (x"40",x"40",x"40",x"40"),
   166 => (x"06",x"7f",x"7f",x"00"),
   167 => (x"7f",x"7f",x"06",x"0c"),
   168 => (x"06",x"7f",x"7f",x"00"),
   169 => (x"7f",x"7f",x"18",x"0c"),
   170 => (x"7f",x"3e",x"00",x"00"),
   171 => (x"3e",x"7f",x"41",x"41"),
   172 => (x"7f",x"7f",x"00",x"00"),
   173 => (x"06",x"0f",x"09",x"09"),
   174 => (x"41",x"7f",x"3e",x"00"),
   175 => (x"40",x"7e",x"7f",x"61"),
   176 => (x"7f",x"7f",x"00",x"00"),
   177 => (x"66",x"7f",x"19",x"09"),
   178 => (x"6f",x"26",x"00",x"00"),
   179 => (x"32",x"7b",x"59",x"4d"),
   180 => (x"01",x"01",x"00",x"00"),
   181 => (x"01",x"01",x"7f",x"7f"),
   182 => (x"7f",x"3f",x"00",x"00"),
   183 => (x"3f",x"7f",x"40",x"40"),
   184 => (x"3f",x"0f",x"00",x"00"),
   185 => (x"0f",x"3f",x"70",x"70"),
   186 => (x"30",x"7f",x"7f",x"00"),
   187 => (x"7f",x"7f",x"30",x"18"),
   188 => (x"36",x"63",x"41",x"00"),
   189 => (x"63",x"36",x"1c",x"1c"),
   190 => (x"06",x"03",x"01",x"41"),
   191 => (x"03",x"06",x"7c",x"7c"),
   192 => (x"59",x"71",x"61",x"01"),
   193 => (x"41",x"43",x"47",x"4d"),
   194 => (x"7f",x"00",x"00",x"00"),
   195 => (x"00",x"41",x"41",x"7f"),
   196 => (x"06",x"03",x"01",x"00"),
   197 => (x"60",x"30",x"18",x"0c"),
   198 => (x"41",x"00",x"00",x"40"),
   199 => (x"00",x"7f",x"7f",x"41"),
   200 => (x"06",x"0c",x"08",x"00"),
   201 => (x"08",x"0c",x"06",x"03"),
   202 => (x"80",x"80",x"80",x"00"),
   203 => (x"80",x"80",x"80",x"80"),
   204 => (x"00",x"00",x"00",x"00"),
   205 => (x"00",x"04",x"07",x"03"),
   206 => (x"74",x"20",x"00",x"00"),
   207 => (x"78",x"7c",x"54",x"54"),
   208 => (x"7f",x"7f",x"00",x"00"),
   209 => (x"38",x"7c",x"44",x"44"),
   210 => (x"7c",x"38",x"00",x"00"),
   211 => (x"00",x"44",x"44",x"44"),
   212 => (x"7c",x"38",x"00",x"00"),
   213 => (x"7f",x"7f",x"44",x"44"),
   214 => (x"7c",x"38",x"00",x"00"),
   215 => (x"18",x"5c",x"54",x"54"),
   216 => (x"7e",x"04",x"00",x"00"),
   217 => (x"00",x"05",x"05",x"7f"),
   218 => (x"bc",x"18",x"00",x"00"),
   219 => (x"7c",x"fc",x"a4",x"a4"),
   220 => (x"7f",x"7f",x"00",x"00"),
   221 => (x"78",x"7c",x"04",x"04"),
   222 => (x"00",x"00",x"00",x"00"),
   223 => (x"00",x"40",x"7d",x"3d"),
   224 => (x"80",x"80",x"00",x"00"),
   225 => (x"00",x"7d",x"fd",x"80"),
   226 => (x"7f",x"7f",x"00",x"00"),
   227 => (x"44",x"6c",x"38",x"10"),
   228 => (x"00",x"00",x"00",x"00"),
   229 => (x"00",x"40",x"7f",x"3f"),
   230 => (x"0c",x"7c",x"7c",x"00"),
   231 => (x"78",x"7c",x"0c",x"18"),
   232 => (x"7c",x"7c",x"00",x"00"),
   233 => (x"78",x"7c",x"04",x"04"),
   234 => (x"7c",x"38",x"00",x"00"),
   235 => (x"38",x"7c",x"44",x"44"),
   236 => (x"fc",x"fc",x"00",x"00"),
   237 => (x"18",x"3c",x"24",x"24"),
   238 => (x"3c",x"18",x"00",x"00"),
   239 => (x"fc",x"fc",x"24",x"24"),
   240 => (x"7c",x"7c",x"00",x"00"),
   241 => (x"08",x"0c",x"04",x"04"),
   242 => (x"5c",x"48",x"00",x"00"),
   243 => (x"20",x"74",x"54",x"54"),
   244 => (x"3f",x"04",x"00",x"00"),
   245 => (x"00",x"44",x"44",x"7f"),
   246 => (x"7c",x"3c",x"00",x"00"),
   247 => (x"7c",x"7c",x"40",x"40"),
   248 => (x"3c",x"1c",x"00",x"00"),
   249 => (x"1c",x"3c",x"60",x"60"),
   250 => (x"60",x"7c",x"3c",x"00"),
   251 => (x"3c",x"7c",x"60",x"30"),
   252 => (x"38",x"6c",x"44",x"00"),
   253 => (x"44",x"6c",x"38",x"10"),
   254 => (x"bc",x"1c",x"00",x"00"),
   255 => (x"1c",x"3c",x"60",x"e0"),
   256 => (x"64",x"44",x"00",x"00"),
   257 => (x"44",x"4c",x"5c",x"74"),
   258 => (x"08",x"08",x"00",x"00"),
   259 => (x"41",x"41",x"77",x"3e"),
   260 => (x"00",x"00",x"00",x"00"),
   261 => (x"00",x"00",x"7f",x"7f"),
   262 => (x"41",x"41",x"00",x"00"),
   263 => (x"08",x"08",x"3e",x"77"),
   264 => (x"01",x"01",x"02",x"00"),
   265 => (x"01",x"02",x"02",x"03"),
   266 => (x"7f",x"7f",x"7f",x"00"),
   267 => (x"7f",x"7f",x"7f",x"7f"),
   268 => (x"1c",x"08",x"08",x"00"),
   269 => (x"7f",x"3e",x"3e",x"1c"),
   270 => (x"3e",x"7f",x"7f",x"7f"),
   271 => (x"08",x"1c",x"1c",x"3e"),
   272 => (x"18",x"10",x"00",x"08"),
   273 => (x"10",x"18",x"7c",x"7c"),
   274 => (x"30",x"10",x"00",x"00"),
   275 => (x"10",x"30",x"7c",x"7c"),
   276 => (x"60",x"30",x"10",x"00"),
   277 => (x"06",x"1e",x"78",x"60"),
   278 => (x"3c",x"66",x"42",x"00"),
   279 => (x"42",x"66",x"3c",x"18"),
   280 => (x"6a",x"38",x"78",x"00"),
   281 => (x"38",x"6c",x"c6",x"c2"),
   282 => (x"00",x"00",x"60",x"00"),
   283 => (x"60",x"00",x"00",x"60"),
   284 => (x"5b",x"5e",x"0e",x"00"),
   285 => (x"1e",x"0e",x"5d",x"5c"),
   286 => (x"f8",x"c2",x"4c",x"71"),
   287 => (x"c0",x"4d",x"bf",x"c9"),
   288 => (x"74",x"1e",x"c0",x"4b"),
   289 => (x"87",x"c7",x"02",x"ab"),
   290 => (x"c0",x"48",x"a6",x"c4"),
   291 => (x"c4",x"87",x"c5",x"78"),
   292 => (x"78",x"c1",x"48",x"a6"),
   293 => (x"73",x"1e",x"66",x"c4"),
   294 => (x"87",x"df",x"ee",x"49"),
   295 => (x"e0",x"c0",x"86",x"c8"),
   296 => (x"87",x"ef",x"ef",x"49"),
   297 => (x"6a",x"4a",x"a5",x"c4"),
   298 => (x"87",x"f0",x"f0",x"49"),
   299 => (x"cb",x"87",x"c6",x"f1"),
   300 => (x"c8",x"83",x"c1",x"85"),
   301 => (x"ff",x"04",x"ab",x"b7"),
   302 => (x"26",x"26",x"87",x"c7"),
   303 => (x"26",x"4c",x"26",x"4d"),
   304 => (x"1e",x"4f",x"26",x"4b"),
   305 => (x"f8",x"c2",x"4a",x"71"),
   306 => (x"f8",x"c2",x"5a",x"cd"),
   307 => (x"78",x"c7",x"48",x"cd"),
   308 => (x"87",x"dd",x"fe",x"49"),
   309 => (x"73",x"1e",x"4f",x"26"),
   310 => (x"c0",x"4a",x"71",x"1e"),
   311 => (x"d3",x"03",x"aa",x"b7"),
   312 => (x"f6",x"e0",x"c2",x"87"),
   313 => (x"87",x"c4",x"05",x"bf"),
   314 => (x"87",x"c2",x"4b",x"c1"),
   315 => (x"e0",x"c2",x"4b",x"c0"),
   316 => (x"87",x"c4",x"5b",x"fa"),
   317 => (x"5a",x"fa",x"e0",x"c2"),
   318 => (x"bf",x"f6",x"e0",x"c2"),
   319 => (x"c1",x"9a",x"c1",x"4a"),
   320 => (x"ec",x"49",x"a2",x"c0"),
   321 => (x"48",x"fc",x"87",x"e8"),
   322 => (x"bf",x"f6",x"e0",x"c2"),
   323 => (x"87",x"ef",x"fe",x"78"),
   324 => (x"c4",x"4a",x"71",x"1e"),
   325 => (x"49",x"72",x"1e",x"66"),
   326 => (x"87",x"dd",x"df",x"ff"),
   327 => (x"1e",x"4f",x"26",x"26"),
   328 => (x"bf",x"f6",x"e0",x"c2"),
   329 => (x"cd",x"dc",x"ff",x"49"),
   330 => (x"c1",x"f8",x"c2",x"87"),
   331 => (x"78",x"bf",x"e8",x"48"),
   332 => (x"48",x"fd",x"f7",x"c2"),
   333 => (x"c2",x"78",x"bf",x"ec"),
   334 => (x"4a",x"bf",x"c1",x"f8"),
   335 => (x"99",x"ff",x"c3",x"49"),
   336 => (x"72",x"2a",x"b7",x"c8"),
   337 => (x"c2",x"b0",x"71",x"48"),
   338 => (x"26",x"58",x"c9",x"f8"),
   339 => (x"5b",x"5e",x"0e",x"4f"),
   340 => (x"71",x"0e",x"5d",x"5c"),
   341 => (x"87",x"c7",x"ff",x"4b"),
   342 => (x"48",x"fc",x"f7",x"c2"),
   343 => (x"49",x"73",x"50",x"c0"),
   344 => (x"87",x"f2",x"db",x"ff"),
   345 => (x"c2",x"4c",x"49",x"70"),
   346 => (x"49",x"ee",x"cb",x"9c"),
   347 => (x"70",x"87",x"cf",x"cb"),
   348 => (x"f7",x"c2",x"4d",x"49"),
   349 => (x"05",x"bf",x"97",x"fc"),
   350 => (x"d0",x"87",x"e4",x"c1"),
   351 => (x"f8",x"c2",x"49",x"66"),
   352 => (x"05",x"99",x"bf",x"c5"),
   353 => (x"66",x"d4",x"87",x"d7"),
   354 => (x"fd",x"f7",x"c2",x"49"),
   355 => (x"cc",x"05",x"99",x"bf"),
   356 => (x"ff",x"49",x"73",x"87"),
   357 => (x"70",x"87",x"ff",x"da"),
   358 => (x"c2",x"c1",x"02",x"98"),
   359 => (x"fd",x"4c",x"c1",x"87"),
   360 => (x"49",x"75",x"87",x"fd"),
   361 => (x"70",x"87",x"e3",x"ca"),
   362 => (x"87",x"c6",x"02",x"98"),
   363 => (x"48",x"fc",x"f7",x"c2"),
   364 => (x"f7",x"c2",x"50",x"c1"),
   365 => (x"05",x"bf",x"97",x"fc"),
   366 => (x"c2",x"87",x"e4",x"c0"),
   367 => (x"49",x"bf",x"c5",x"f8"),
   368 => (x"05",x"99",x"66",x"d0"),
   369 => (x"c2",x"87",x"d6",x"ff"),
   370 => (x"49",x"bf",x"fd",x"f7"),
   371 => (x"05",x"99",x"66",x"d4"),
   372 => (x"73",x"87",x"ca",x"ff"),
   373 => (x"fd",x"d9",x"ff",x"49"),
   374 => (x"05",x"98",x"70",x"87"),
   375 => (x"74",x"87",x"fe",x"fe"),
   376 => (x"87",x"d7",x"fb",x"48"),
   377 => (x"5c",x"5b",x"5e",x"0e"),
   378 => (x"86",x"f4",x"0e",x"5d"),
   379 => (x"ec",x"4c",x"4d",x"c0"),
   380 => (x"a6",x"c4",x"7e",x"bf"),
   381 => (x"c9",x"f8",x"c2",x"48"),
   382 => (x"1e",x"c1",x"78",x"bf"),
   383 => (x"49",x"c7",x"1e",x"c0"),
   384 => (x"c8",x"87",x"ca",x"fd"),
   385 => (x"02",x"98",x"70",x"86"),
   386 => (x"49",x"ff",x"87",x"ce"),
   387 => (x"c1",x"87",x"c7",x"fb"),
   388 => (x"d9",x"ff",x"49",x"da"),
   389 => (x"4d",x"c1",x"87",x"c0"),
   390 => (x"97",x"fc",x"f7",x"c2"),
   391 => (x"87",x"c3",x"02",x"bf"),
   392 => (x"c2",x"87",x"c0",x"c9"),
   393 => (x"4b",x"bf",x"c1",x"f8"),
   394 => (x"bf",x"f6",x"e0",x"c2"),
   395 => (x"87",x"eb",x"c0",x"05"),
   396 => (x"ff",x"49",x"fd",x"c3"),
   397 => (x"c3",x"87",x"df",x"d8"),
   398 => (x"d8",x"ff",x"49",x"fa"),
   399 => (x"49",x"73",x"87",x"d8"),
   400 => (x"71",x"99",x"ff",x"c3"),
   401 => (x"fb",x"49",x"c0",x"1e"),
   402 => (x"49",x"73",x"87",x"c6"),
   403 => (x"71",x"29",x"b7",x"c8"),
   404 => (x"fa",x"49",x"c1",x"1e"),
   405 => (x"86",x"c8",x"87",x"fa"),
   406 => (x"c2",x"87",x"c1",x"c6"),
   407 => (x"4b",x"bf",x"c5",x"f8"),
   408 => (x"87",x"dd",x"02",x"9b"),
   409 => (x"bf",x"f2",x"e0",x"c2"),
   410 => (x"87",x"de",x"c7",x"49"),
   411 => (x"c4",x"05",x"98",x"70"),
   412 => (x"d2",x"4b",x"c0",x"87"),
   413 => (x"49",x"e0",x"c2",x"87"),
   414 => (x"c2",x"87",x"c3",x"c7"),
   415 => (x"c6",x"58",x"f6",x"e0"),
   416 => (x"f2",x"e0",x"c2",x"87"),
   417 => (x"73",x"78",x"c0",x"48"),
   418 => (x"05",x"99",x"c2",x"49"),
   419 => (x"eb",x"c3",x"87",x"ce"),
   420 => (x"c1",x"d7",x"ff",x"49"),
   421 => (x"c2",x"49",x"70",x"87"),
   422 => (x"87",x"c2",x"02",x"99"),
   423 => (x"49",x"73",x"4c",x"fb"),
   424 => (x"ce",x"05",x"99",x"c1"),
   425 => (x"49",x"f4",x"c3",x"87"),
   426 => (x"87",x"ea",x"d6",x"ff"),
   427 => (x"99",x"c2",x"49",x"70"),
   428 => (x"fa",x"87",x"c2",x"02"),
   429 => (x"c8",x"49",x"73",x"4c"),
   430 => (x"87",x"ce",x"05",x"99"),
   431 => (x"ff",x"49",x"f5",x"c3"),
   432 => (x"70",x"87",x"d3",x"d6"),
   433 => (x"02",x"99",x"c2",x"49"),
   434 => (x"f8",x"c2",x"87",x"d5"),
   435 => (x"ca",x"02",x"bf",x"cd"),
   436 => (x"88",x"c1",x"48",x"87"),
   437 => (x"58",x"d1",x"f8",x"c2"),
   438 => (x"ff",x"87",x"c2",x"c0"),
   439 => (x"73",x"4d",x"c1",x"4c"),
   440 => (x"05",x"99",x"c4",x"49"),
   441 => (x"f2",x"c3",x"87",x"ce"),
   442 => (x"e9",x"d5",x"ff",x"49"),
   443 => (x"c2",x"49",x"70",x"87"),
   444 => (x"87",x"dc",x"02",x"99"),
   445 => (x"bf",x"cd",x"f8",x"c2"),
   446 => (x"b7",x"c7",x"48",x"7e"),
   447 => (x"cb",x"c0",x"03",x"a8"),
   448 => (x"c1",x"48",x"6e",x"87"),
   449 => (x"d1",x"f8",x"c2",x"80"),
   450 => (x"87",x"c2",x"c0",x"58"),
   451 => (x"4d",x"c1",x"4c",x"fe"),
   452 => (x"ff",x"49",x"fd",x"c3"),
   453 => (x"70",x"87",x"ff",x"d4"),
   454 => (x"02",x"99",x"c2",x"49"),
   455 => (x"c2",x"87",x"d5",x"c0"),
   456 => (x"02",x"bf",x"cd",x"f8"),
   457 => (x"c2",x"87",x"c9",x"c0"),
   458 => (x"c0",x"48",x"cd",x"f8"),
   459 => (x"87",x"c2",x"c0",x"78"),
   460 => (x"4d",x"c1",x"4c",x"fd"),
   461 => (x"ff",x"49",x"fa",x"c3"),
   462 => (x"70",x"87",x"db",x"d4"),
   463 => (x"02",x"99",x"c2",x"49"),
   464 => (x"c2",x"87",x"d9",x"c0"),
   465 => (x"48",x"bf",x"cd",x"f8"),
   466 => (x"03",x"a8",x"b7",x"c7"),
   467 => (x"c2",x"87",x"c9",x"c0"),
   468 => (x"c7",x"48",x"cd",x"f8"),
   469 => (x"87",x"c2",x"c0",x"78"),
   470 => (x"4d",x"c1",x"4c",x"fc"),
   471 => (x"03",x"ac",x"b7",x"c0"),
   472 => (x"c4",x"87",x"d1",x"c0"),
   473 => (x"d8",x"c1",x"4a",x"66"),
   474 => (x"c0",x"02",x"6a",x"82"),
   475 => (x"4b",x"6a",x"87",x"c6"),
   476 => (x"0f",x"73",x"49",x"74"),
   477 => (x"f0",x"c3",x"1e",x"c0"),
   478 => (x"49",x"da",x"c1",x"1e"),
   479 => (x"c8",x"87",x"ce",x"f7"),
   480 => (x"02",x"98",x"70",x"86"),
   481 => (x"c8",x"87",x"e2",x"c0"),
   482 => (x"f8",x"c2",x"48",x"a6"),
   483 => (x"c8",x"78",x"bf",x"cd"),
   484 => (x"91",x"cb",x"49",x"66"),
   485 => (x"71",x"48",x"66",x"c4"),
   486 => (x"6e",x"7e",x"70",x"80"),
   487 => (x"c8",x"c0",x"02",x"bf"),
   488 => (x"4b",x"bf",x"6e",x"87"),
   489 => (x"73",x"49",x"66",x"c8"),
   490 => (x"02",x"9d",x"75",x"0f"),
   491 => (x"c2",x"87",x"c8",x"c0"),
   492 => (x"49",x"bf",x"cd",x"f8"),
   493 => (x"c2",x"87",x"fa",x"f2"),
   494 => (x"02",x"bf",x"fa",x"e0"),
   495 => (x"49",x"87",x"dd",x"c0"),
   496 => (x"70",x"87",x"c7",x"c2"),
   497 => (x"d3",x"c0",x"02",x"98"),
   498 => (x"cd",x"f8",x"c2",x"87"),
   499 => (x"e0",x"f2",x"49",x"bf"),
   500 => (x"f4",x"49",x"c0",x"87"),
   501 => (x"e0",x"c2",x"87",x"c0"),
   502 => (x"78",x"c0",x"48",x"fa"),
   503 => (x"da",x"f3",x"8e",x"f4"),
   504 => (x"5b",x"5e",x"0e",x"87"),
   505 => (x"1e",x"0e",x"5d",x"5c"),
   506 => (x"f8",x"c2",x"4c",x"71"),
   507 => (x"c1",x"49",x"bf",x"c9"),
   508 => (x"c1",x"4d",x"a1",x"cd"),
   509 => (x"7e",x"69",x"81",x"d1"),
   510 => (x"cf",x"02",x"9c",x"74"),
   511 => (x"4b",x"a5",x"c4",x"87"),
   512 => (x"f8",x"c2",x"7b",x"74"),
   513 => (x"f2",x"49",x"bf",x"c9"),
   514 => (x"7b",x"6e",x"87",x"f9"),
   515 => (x"c4",x"05",x"9c",x"74"),
   516 => (x"c2",x"4b",x"c0",x"87"),
   517 => (x"73",x"4b",x"c1",x"87"),
   518 => (x"87",x"fa",x"f2",x"49"),
   519 => (x"c7",x"02",x"66",x"d4"),
   520 => (x"87",x"da",x"49",x"87"),
   521 => (x"87",x"c2",x"4a",x"70"),
   522 => (x"e0",x"c2",x"4a",x"c0"),
   523 => (x"f2",x"26",x"5a",x"fe"),
   524 => (x"00",x"00",x"87",x"c9"),
   525 => (x"00",x"00",x"00",x"00"),
   526 => (x"00",x"00",x"00",x"00"),
   527 => (x"71",x"1e",x"00",x"00"),
   528 => (x"bf",x"c8",x"ff",x"4a"),
   529 => (x"48",x"a1",x"72",x"49"),
   530 => (x"ff",x"1e",x"4f",x"26"),
   531 => (x"fe",x"89",x"bf",x"c8"),
   532 => (x"c0",x"c0",x"c0",x"c0"),
   533 => (x"c4",x"01",x"a9",x"c0"),
   534 => (x"c2",x"4a",x"c0",x"87"),
   535 => (x"72",x"4a",x"c1",x"87"),
   536 => (x"1e",x"4f",x"26",x"48"),
   537 => (x"bf",x"f1",x"e2",x"c2"),
   538 => (x"c2",x"b9",x"c1",x"49"),
   539 => (x"ff",x"59",x"f5",x"e2"),
   540 => (x"ff",x"c3",x"48",x"d4"),
   541 => (x"48",x"d0",x"ff",x"78"),
   542 => (x"ff",x"78",x"e1",x"c0"),
   543 => (x"78",x"c1",x"48",x"d4"),
   544 => (x"78",x"71",x"31",x"c4"),
   545 => (x"c0",x"48",x"d0",x"ff"),
   546 => (x"4f",x"26",x"78",x"e0"),
   547 => (x"e5",x"e2",x"c2",x"1e"),
   548 => (x"f0",x"f2",x"c2",x"1e"),
   549 => (x"f9",x"fb",x"fd",x"49"),
   550 => (x"70",x"86",x"c4",x"87"),
   551 => (x"87",x"c3",x"02",x"98"),
   552 => (x"26",x"87",x"c0",x"ff"),
   553 => (x"4b",x"35",x"31",x"4f"),
   554 => (x"20",x"20",x"5a",x"48"),
   555 => (x"47",x"46",x"43",x"20"),
   556 => (x"00",x"00",x"00",x"00"),
   557 => (x"5b",x"5e",x"0e",x"00"),
   558 => (x"c2",x"0e",x"5d",x"5c"),
   559 => (x"4a",x"bf",x"fd",x"f7"),
   560 => (x"bf",x"de",x"e4",x"c2"),
   561 => (x"bc",x"72",x"4c",x"49"),
   562 => (x"c6",x"ff",x"4d",x"71"),
   563 => (x"4b",x"c0",x"87",x"df"),
   564 => (x"99",x"d0",x"49",x"74"),
   565 => (x"87",x"e7",x"c0",x"02"),
   566 => (x"c8",x"48",x"d0",x"ff"),
   567 => (x"d4",x"ff",x"78",x"e1"),
   568 => (x"75",x"78",x"c5",x"48"),
   569 => (x"02",x"99",x"d0",x"49"),
   570 => (x"f0",x"c3",x"87",x"c3"),
   571 => (x"cc",x"e5",x"c2",x"78"),
   572 => (x"11",x"81",x"73",x"49"),
   573 => (x"08",x"d4",x"ff",x"48"),
   574 => (x"48",x"d0",x"ff",x"78"),
   575 => (x"c1",x"78",x"e0",x"c0"),
   576 => (x"c8",x"83",x"2d",x"2c"),
   577 => (x"c7",x"ff",x"04",x"ab"),
   578 => (x"d8",x"c5",x"ff",x"87"),
   579 => (x"de",x"e4",x"c2",x"87"),
   580 => (x"fd",x"f7",x"c2",x"48"),
   581 => (x"4d",x"26",x"78",x"bf"),
   582 => (x"4b",x"26",x"4c",x"26"),
   583 => (x"00",x"00",x"4f",x"26"),
   584 => (x"c1",x"1e",x"00",x"00"),
   585 => (x"de",x"48",x"d0",x"e7"),
   586 => (x"f5",x"e4",x"c2",x"50"),
   587 => (x"e2",x"d9",x"fe",x"49"),
   588 => (x"26",x"48",x"c0",x"87"),
   589 => (x"4f",x"54",x"4a",x"4f"),
   590 => (x"55",x"52",x"54",x"55"),
   591 => (x"43",x"52",x"41",x"4e"),
   592 => (x"df",x"f2",x"1e",x"00"),
   593 => (x"87",x"ed",x"fd",x"87"),
   594 => (x"4f",x"26",x"87",x"f8"),
   595 => (x"25",x"26",x"1e",x"16"),
   596 => (x"3e",x"3d",x"36",x"2e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

