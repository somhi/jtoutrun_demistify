library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c0f8c287",
    12 => x"86c0c84e",
    13 => x"49c0f8c2",
    14 => x"48c0e5c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087ede5",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"8148731e",
    47 => x"7205a973",
    48 => x"2687f953",
    49 => x"4a711e4f",
    50 => x"484966c4",
    51 => x"a6c888c1",
    52 => x"02997158",
    53 => x"d4ff87d6",
    54 => x"78ffc348",
    55 => x"66c45268",
    56 => x"88c14849",
    57 => x"7158a6c8",
    58 => x"87ea0599",
    59 => x"731e4f26",
    60 => x"4bd4ff1e",
    61 => x"6b7bffc3",
    62 => x"7bffc34a",
    63 => x"32c8496b",
    64 => x"ffc3b172",
    65 => x"c84a6b7b",
    66 => x"c3b27131",
    67 => x"496b7bff",
    68 => x"b17232c8",
    69 => x"87c44871",
    70 => x"4c264d26",
    71 => x"4f264b26",
    72 => x"5c5b5e0e",
    73 => x"4a710e5d",
    74 => x"724cd4ff",
    75 => x"99ffc349",
    76 => x"e5c27c71",
    77 => x"c805bfc0",
    78 => x"4866d087",
    79 => x"a6d430c9",
    80 => x"4966d058",
    81 => x"ffc329d8",
    82 => x"d07c7199",
    83 => x"29d04966",
    84 => x"7199ffc3",
    85 => x"4966d07c",
    86 => x"ffc329c8",
    87 => x"d07c7199",
    88 => x"ffc34966",
    89 => x"727c7199",
    90 => x"c329d049",
    91 => x"7c7199ff",
    92 => x"f0c94b6c",
    93 => x"ffc34dff",
    94 => x"87d005ab",
    95 => x"6c7cffc3",
    96 => x"028dc14b",
    97 => x"ffc387c6",
    98 => x"87f002ab",
    99 => x"c7fe4873",
   100 => x"49c01e87",
   101 => x"c348d4ff",
   102 => x"81c178ff",
   103 => x"a9b7c8c3",
   104 => x"2687f104",
   105 => x"1e731e4f",
   106 => x"f8c487e7",
   107 => x"1ec04bdf",
   108 => x"c1f0ffc0",
   109 => x"e7fd49f7",
   110 => x"c186c487",
   111 => x"eac005a8",
   112 => x"48d4ff87",
   113 => x"c178ffc3",
   114 => x"c0c0c0c0",
   115 => x"e1c01ec0",
   116 => x"49e9c1f0",
   117 => x"c487c9fd",
   118 => x"05987086",
   119 => x"d4ff87ca",
   120 => x"78ffc348",
   121 => x"87cb48c1",
   122 => x"c187e6fe",
   123 => x"fdfe058b",
   124 => x"fc48c087",
   125 => x"731e87e6",
   126 => x"48d4ff1e",
   127 => x"d378ffc3",
   128 => x"c01ec04b",
   129 => x"c1c1f0ff",
   130 => x"87d4fc49",
   131 => x"987086c4",
   132 => x"ff87ca05",
   133 => x"ffc348d4",
   134 => x"cb48c178",
   135 => x"87f1fd87",
   136 => x"ff058bc1",
   137 => x"48c087db",
   138 => x"0e87f1fb",
   139 => x"0e5c5b5e",
   140 => x"fd4cd4ff",
   141 => x"eac687db",
   142 => x"f0e1c01e",
   143 => x"fb49c8c1",
   144 => x"86c487de",
   145 => x"c802a8c1",
   146 => x"87eafe87",
   147 => x"e2c148c0",
   148 => x"87dafa87",
   149 => x"ffcf4970",
   150 => x"eac699ff",
   151 => x"87c802a9",
   152 => x"c087d3fe",
   153 => x"87cbc148",
   154 => x"c07cffc3",
   155 => x"f4fc4bf1",
   156 => x"02987087",
   157 => x"c087ebc0",
   158 => x"f0ffc01e",
   159 => x"fa49fac1",
   160 => x"86c487de",
   161 => x"d9059870",
   162 => x"7cffc387",
   163 => x"ffc3496c",
   164 => x"7c7c7c7c",
   165 => x"0299c0c1",
   166 => x"48c187c4",
   167 => x"48c087d5",
   168 => x"abc287d1",
   169 => x"c087c405",
   170 => x"c187c848",
   171 => x"fdfe058b",
   172 => x"f948c087",
   173 => x"731e87e4",
   174 => x"c0e5c21e",
   175 => x"c778c148",
   176 => x"48d0ff4b",
   177 => x"c8fb78c2",
   178 => x"48d0ff87",
   179 => x"1ec078c3",
   180 => x"c1d0e5c0",
   181 => x"c7f949c0",
   182 => x"c186c487",
   183 => x"87c105a8",
   184 => x"05abc24b",
   185 => x"48c087c5",
   186 => x"c187f9c0",
   187 => x"d0ff058b",
   188 => x"87f7fc87",
   189 => x"58c4e5c2",
   190 => x"cd059870",
   191 => x"c01ec187",
   192 => x"d0c1f0ff",
   193 => x"87d8f849",
   194 => x"d4ff86c4",
   195 => x"78ffc348",
   196 => x"c287fcc2",
   197 => x"ff58c8e5",
   198 => x"78c248d0",
   199 => x"c348d4ff",
   200 => x"48c178ff",
   201 => x"0e87f5f7",
   202 => x"5d5c5b5e",
   203 => x"c04b710e",
   204 => x"cdeec54c",
   205 => x"d4ff4adf",
   206 => x"78ffc348",
   207 => x"fec34968",
   208 => x"fdc005a9",
   209 => x"734d7087",
   210 => x"87cc029b",
   211 => x"731e66d0",
   212 => x"87f1f549",
   213 => x"87d686c4",
   214 => x"c448d0ff",
   215 => x"ffc378d1",
   216 => x"4866d07d",
   217 => x"a6d488c1",
   218 => x"05987058",
   219 => x"d4ff87f0",
   220 => x"78ffc348",
   221 => x"059b7378",
   222 => x"d0ff87c5",
   223 => x"c178d048",
   224 => x"8ac14c4a",
   225 => x"87eefe05",
   226 => x"cbf64874",
   227 => x"1e731e87",
   228 => x"4bc04a71",
   229 => x"c348d4ff",
   230 => x"d0ff78ff",
   231 => x"78c3c448",
   232 => x"c348d4ff",
   233 => x"1e7278ff",
   234 => x"c1f0ffc0",
   235 => x"eff549d1",
   236 => x"7086c487",
   237 => x"87d20598",
   238 => x"cc1ec0c8",
   239 => x"e6fd4966",
   240 => x"7086c487",
   241 => x"48d0ff4b",
   242 => x"487378c2",
   243 => x"0e87cdf5",
   244 => x"5d5c5b5e",
   245 => x"c01ec00e",
   246 => x"c9c1f0ff",
   247 => x"87c0f549",
   248 => x"e5c21ed2",
   249 => x"fefc49c8",
   250 => x"c086c887",
   251 => x"d284c14c",
   252 => x"f804acb7",
   253 => x"c8e5c287",
   254 => x"c349bf97",
   255 => x"c0c199c0",
   256 => x"e7c005a9",
   257 => x"cfe5c287",
   258 => x"d049bf97",
   259 => x"d0e5c231",
   260 => x"c84abf97",
   261 => x"c2b17232",
   262 => x"bf97d1e5",
   263 => x"4c71b14a",
   264 => x"ffffffcf",
   265 => x"ca84c19c",
   266 => x"87e7c134",
   267 => x"97d1e5c2",
   268 => x"31c149bf",
   269 => x"e5c299c6",
   270 => x"4abf97d2",
   271 => x"722ab7c7",
   272 => x"cde5c2b1",
   273 => x"4d4abf97",
   274 => x"e5c29dcf",
   275 => x"4abf97ce",
   276 => x"32ca9ac3",
   277 => x"97cfe5c2",
   278 => x"33c24bbf",
   279 => x"e5c2b273",
   280 => x"4bbf97d0",
   281 => x"c69bc0c3",
   282 => x"b2732bb7",
   283 => x"48c181c2",
   284 => x"49703071",
   285 => x"307548c1",
   286 => x"4c724d70",
   287 => x"947184c1",
   288 => x"adb7c0c8",
   289 => x"c187cc06",
   290 => x"c82db734",
   291 => x"01adb7c0",
   292 => x"7487f4ff",
   293 => x"87c0f248",
   294 => x"5c5b5e0e",
   295 => x"86f80e5d",
   296 => x"48eeedc2",
   297 => x"e5c278c0",
   298 => x"49c01ee6",
   299 => x"c487defb",
   300 => x"05987086",
   301 => x"48c087c5",
   302 => x"c087cec9",
   303 => x"c07ec14d",
   304 => x"49bfd8f5",
   305 => x"4adce6c2",
   306 => x"ee4bc871",
   307 => x"987087dc",
   308 => x"c087c205",
   309 => x"d4f5c07e",
   310 => x"e6c249bf",
   311 => x"c8714af8",
   312 => x"87c6ee4b",
   313 => x"c2059870",
   314 => x"6e7ec087",
   315 => x"87fdc002",
   316 => x"bfececc2",
   317 => x"e4edc24d",
   318 => x"487ebf9f",
   319 => x"a8ead6c5",
   320 => x"c287c705",
   321 => x"4dbfecec",
   322 => x"486e87ce",
   323 => x"a8d5e9ca",
   324 => x"c087c502",
   325 => x"87f1c748",
   326 => x"1ee6e5c2",
   327 => x"ecf94975",
   328 => x"7086c487",
   329 => x"87c50598",
   330 => x"dcc748c0",
   331 => x"d4f5c087",
   332 => x"e6c249bf",
   333 => x"c8714af8",
   334 => x"87eeec4b",
   335 => x"c8059870",
   336 => x"eeedc287",
   337 => x"da78c148",
   338 => x"d8f5c087",
   339 => x"e6c249bf",
   340 => x"c8714adc",
   341 => x"87d2ec4b",
   342 => x"c0029870",
   343 => x"48c087c5",
   344 => x"c287e6c6",
   345 => x"bf97e4ed",
   346 => x"a9d5c149",
   347 => x"87cdc005",
   348 => x"97e5edc2",
   349 => x"eac249bf",
   350 => x"c5c002a9",
   351 => x"c648c087",
   352 => x"e5c287c7",
   353 => x"7ebf97e6",
   354 => x"a8e9c348",
   355 => x"87cec002",
   356 => x"ebc3486e",
   357 => x"c5c002a8",
   358 => x"c548c087",
   359 => x"e5c287eb",
   360 => x"49bf97f1",
   361 => x"ccc00599",
   362 => x"f2e5c287",
   363 => x"c249bf97",
   364 => x"c5c002a9",
   365 => x"c548c087",
   366 => x"e5c287cf",
   367 => x"48bf97f3",
   368 => x"58eaedc2",
   369 => x"c1484c70",
   370 => x"eeedc288",
   371 => x"f4e5c258",
   372 => x"7549bf97",
   373 => x"f5e5c281",
   374 => x"c84abf97",
   375 => x"7ea17232",
   376 => x"48fbf1c2",
   377 => x"e5c2786e",
   378 => x"48bf97f6",
   379 => x"c258a6c8",
   380 => x"02bfeeed",
   381 => x"c087d4c2",
   382 => x"49bfd4f5",
   383 => x"4af8e6c2",
   384 => x"e94bc871",
   385 => x"987087e4",
   386 => x"87c5c002",
   387 => x"f8c348c0",
   388 => x"e6edc287",
   389 => x"f2c24cbf",
   390 => x"e6c25ccf",
   391 => x"49bf97cb",
   392 => x"e6c231c8",
   393 => x"4abf97ca",
   394 => x"e6c249a1",
   395 => x"4abf97cc",
   396 => x"a17232d0",
   397 => x"cde6c249",
   398 => x"d84abf97",
   399 => x"49a17232",
   400 => x"c29166c4",
   401 => x"81bffbf1",
   402 => x"59c3f2c2",
   403 => x"97d3e6c2",
   404 => x"32c84abf",
   405 => x"97d2e6c2",
   406 => x"4aa24bbf",
   407 => x"97d4e6c2",
   408 => x"33d04bbf",
   409 => x"c24aa273",
   410 => x"bf97d5e6",
   411 => x"d89bcf4b",
   412 => x"4aa27333",
   413 => x"5ac7f2c2",
   414 => x"bfc3f2c2",
   415 => x"748ac24a",
   416 => x"c7f2c292",
   417 => x"78a17248",
   418 => x"c287cac1",
   419 => x"bf97f8e5",
   420 => x"c231c849",
   421 => x"bf97f7e5",
   422 => x"c249a14a",
   423 => x"c259f6ed",
   424 => x"49bff2ed",
   425 => x"ffc731c5",
   426 => x"c229c981",
   427 => x"c259cff2",
   428 => x"bf97fde5",
   429 => x"c232c84a",
   430 => x"bf97fce5",
   431 => x"c44aa24b",
   432 => x"826e9266",
   433 => x"5acbf2c2",
   434 => x"48c3f2c2",
   435 => x"f1c278c0",
   436 => x"a17248ff",
   437 => x"cff2c278",
   438 => x"c3f2c248",
   439 => x"f2c278bf",
   440 => x"f2c248d3",
   441 => x"c278bfc7",
   442 => x"02bfeeed",
   443 => x"7487c9c0",
   444 => x"7030c448",
   445 => x"87c9c07e",
   446 => x"bfcbf2c2",
   447 => x"7030c448",
   448 => x"f2edc27e",
   449 => x"c1786e48",
   450 => x"268ef848",
   451 => x"264c264d",
   452 => x"0e4f264b",
   453 => x"5d5c5b5e",
   454 => x"c24a710e",
   455 => x"02bfeeed",
   456 => x"4b7287cb",
   457 => x"4c722bc7",
   458 => x"c99cffc1",
   459 => x"c84b7287",
   460 => x"c34c722b",
   461 => x"f1c29cff",
   462 => x"c083bffb",
   463 => x"abbfd0f5",
   464 => x"c087d902",
   465 => x"c25bd4f5",
   466 => x"731ee6e5",
   467 => x"87fdf049",
   468 => x"987086c4",
   469 => x"c087c505",
   470 => x"87e6c048",
   471 => x"bfeeedc2",
   472 => x"7487d202",
   473 => x"c291c449",
   474 => x"6981e6e5",
   475 => x"ffffcf4d",
   476 => x"cb9dffff",
   477 => x"c2497487",
   478 => x"e6e5c291",
   479 => x"4d699f81",
   480 => x"c6fe4875",
   481 => x"5b5e0e87",
   482 => x"f80e5d5c",
   483 => x"9c4c7186",
   484 => x"c087c505",
   485 => x"87c1c348",
   486 => x"6e7ea4c8",
   487 => x"d878c048",
   488 => x"87c70266",
   489 => x"bf9766d8",
   490 => x"c087c505",
   491 => x"87e9c248",
   492 => x"49c11ec0",
   493 => x"c487fdce",
   494 => x"9d4d7086",
   495 => x"87c2c102",
   496 => x"4af6edc2",
   497 => x"e24966d8",
   498 => x"987087c5",
   499 => x"87f2c002",
   500 => x"66d84a75",
   501 => x"e24bcb49",
   502 => x"987087ea",
   503 => x"87e2c002",
   504 => x"9d751ec0",
   505 => x"c887c702",
   506 => x"78c048a6",
   507 => x"a6c887c5",
   508 => x"c878c148",
   509 => x"fbcd4966",
   510 => x"7086c487",
   511 => x"fe059d4d",
   512 => x"9d7587fe",
   513 => x"87cfc102",
   514 => x"6e49a5dc",
   515 => x"da786948",
   516 => x"a6c449a5",
   517 => x"78a4c448",
   518 => x"c448699f",
   519 => x"c2780866",
   520 => x"02bfeeed",
   521 => x"a5d487d2",
   522 => x"49699f49",
   523 => x"99ffffc0",
   524 => x"30d04871",
   525 => x"87c27e70",
   526 => x"496e7ec0",
   527 => x"bf66c448",
   528 => x"0866c480",
   529 => x"cc7cc078",
   530 => x"66c449a4",
   531 => x"a4d079bf",
   532 => x"c179c049",
   533 => x"c087c248",
   534 => x"fa8ef848",
   535 => x"5e0e87ed",
   536 => x"0e5d5c5b",
   537 => x"029c4c71",
   538 => x"c887cac1",
   539 => x"026949a4",
   540 => x"d087c2c1",
   541 => x"496c4a66",
   542 => x"5aa6d482",
   543 => x"b94d66d0",
   544 => x"bfeaedc2",
   545 => x"72baff4a",
   546 => x"02997199",
   547 => x"c487e4c0",
   548 => x"496b4ba4",
   549 => x"7087fcf9",
   550 => x"e6edc27b",
   551 => x"816c49bf",
   552 => x"b9757c71",
   553 => x"bfeaedc2",
   554 => x"72baff4a",
   555 => x"05997199",
   556 => x"7587dcff",
   557 => x"87d3f97c",
   558 => x"711e731e",
   559 => x"c7029b4b",
   560 => x"49a3c887",
   561 => x"87c50569",
   562 => x"f7c048c0",
   563 => x"fff1c287",
   564 => x"a3c44abf",
   565 => x"c2496949",
   566 => x"e6edc289",
   567 => x"a27191bf",
   568 => x"eaedc24a",
   569 => x"996b49bf",
   570 => x"c04aa271",
   571 => x"c85ad4f5",
   572 => x"49721e66",
   573 => x"c487d6ea",
   574 => x"05987086",
   575 => x"48c087c4",
   576 => x"48c187c2",
   577 => x"0e87c8f8",
   578 => x"0e5c5b5e",
   579 => x"d04b711e",
   580 => x"2cc94c66",
   581 => x"c1029b73",
   582 => x"a3c887d4",
   583 => x"c1026949",
   584 => x"edc287cc",
   585 => x"ff49bfea",
   586 => x"994a6bb9",
   587 => x"03ac717e",
   588 => x"7bc087d1",
   589 => x"c049a3d0",
   590 => x"4aa3cc79",
   591 => x"6a49a3c4",
   592 => x"7287c279",
   593 => x"029c748c",
   594 => x"4987e3c0",
   595 => x"fc49731e",
   596 => x"86c487cc",
   597 => x"c74966d0",
   598 => x"cb0299ff",
   599 => x"e6e5c287",
   600 => x"fd49731e",
   601 => x"86c487d2",
   602 => x"d049a3d0",
   603 => x"f6267966",
   604 => x"5e0e87db",
   605 => x"0e5d5c5b",
   606 => x"a6d086f0",
   607 => x"66e4c059",
   608 => x"0266cc4b",
   609 => x"c84887ca",
   610 => x"6e7e7080",
   611 => x"87c505bf",
   612 => x"ecc348c0",
   613 => x"4c66cc87",
   614 => x"497384d0",
   615 => x"6c48a6c4",
   616 => x"8166c478",
   617 => x"bf6e80c4",
   618 => x"a966c878",
   619 => x"4987c606",
   620 => x"718966c4",
   621 => x"abb7c04b",
   622 => x"4887c401",
   623 => x"c487c2c3",
   624 => x"ffc74866",
   625 => x"6e7e7098",
   626 => x"87c9c102",
   627 => x"6e49c0c8",
   628 => x"c24a7189",
   629 => x"6e4de6e5",
   630 => x"aab77385",
   631 => x"4a87c106",
   632 => x"c4484972",
   633 => x"7c708066",
   634 => x"c1498b72",
   635 => x"0299718a",
   636 => x"e0c087d9",
   637 => x"50154866",
   638 => x"4866e0c0",
   639 => x"e4c080c1",
   640 => x"497258a6",
   641 => x"99718ac1",
   642 => x"c187e705",
   643 => x"4966d01e",
   644 => x"c487cbf9",
   645 => x"abb7c086",
   646 => x"87e3c106",
   647 => x"4d66e0c0",
   648 => x"abb7ffc7",
   649 => x"87e2c006",
   650 => x"66d01e75",
   651 => x"87c8fa49",
   652 => x"6c85c0c8",
   653 => x"80c0c848",
   654 => x"c0c87c70",
   655 => x"d41ec18b",
   656 => x"d9f84966",
   657 => x"c086c887",
   658 => x"e5c287ee",
   659 => x"66d01ee6",
   660 => x"87e4f949",
   661 => x"e5c286c4",
   662 => x"49734ae6",
   663 => x"70806c48",
   664 => x"c149737c",
   665 => x"0299718b",
   666 => x"971287ce",
   667 => x"7385c17d",
   668 => x"718bc149",
   669 => x"87f20599",
   670 => x"01abb7c0",
   671 => x"c187e1fe",
   672 => x"f28ef048",
   673 => x"5e0e87c5",
   674 => x"0e5d5c5b",
   675 => x"029b4b71",
   676 => x"a3c887c7",
   677 => x"c5056d4d",
   678 => x"c048ff87",
   679 => x"a3d087fd",
   680 => x"c7496c4c",
   681 => x"d80599ff",
   682 => x"c9026c87",
   683 => x"731ec187",
   684 => x"87eaf649",
   685 => x"e5c286c4",
   686 => x"49731ee6",
   687 => x"c487f9f7",
   688 => x"6d4a6c86",
   689 => x"87c404aa",
   690 => x"87cf48ff",
   691 => x"727ca2c1",
   692 => x"99ffc749",
   693 => x"81e6e5c2",
   694 => x"f0486997",
   695 => x"731e87ed",
   696 => x"9b4b711e",
   697 => x"87e4c002",
   698 => x"5bd3f2c2",
   699 => x"8ac24a73",
   700 => x"bfe6edc2",
   701 => x"f1c29249",
   702 => x"7248bfff",
   703 => x"d7f2c280",
   704 => x"c4487158",
   705 => x"f6edc230",
   706 => x"87edc058",
   707 => x"48cff2c2",
   708 => x"bfc3f2c2",
   709 => x"d3f2c278",
   710 => x"c7f2c248",
   711 => x"edc278bf",
   712 => x"c902bfee",
   713 => x"e6edc287",
   714 => x"31c449bf",
   715 => x"f2c287c7",
   716 => x"c449bfcb",
   717 => x"f6edc231",
   718 => x"87d3ef59",
   719 => x"5c5b5e0e",
   720 => x"c04a710e",
   721 => x"029a724b",
   722 => x"da87e1c0",
   723 => x"699f49a2",
   724 => x"eeedc24b",
   725 => x"87cf02bf",
   726 => x"9f49a2d4",
   727 => x"c04c4969",
   728 => x"d09cffff",
   729 => x"c087c234",
   730 => x"b349744c",
   731 => x"edfd4973",
   732 => x"87d9ee87",
   733 => x"5c5b5e0e",
   734 => x"86f40e5d",
   735 => x"7ec04a71",
   736 => x"d8029a72",
   737 => x"e2e5c287",
   738 => x"c278c048",
   739 => x"c248dae5",
   740 => x"78bfd3f2",
   741 => x"48dee5c2",
   742 => x"bfcff2c2",
   743 => x"c3eec278",
   744 => x"c250c048",
   745 => x"49bff2ed",
   746 => x"bfe2e5c2",
   747 => x"03aa714a",
   748 => x"7287cac4",
   749 => x"0599cf49",
   750 => x"c087eac0",
   751 => x"c248d0f5",
   752 => x"78bfdae5",
   753 => x"1ee6e5c2",
   754 => x"bfdae5c2",
   755 => x"dae5c249",
   756 => x"78a1c148",
   757 => x"f4deff71",
   758 => x"c086c487",
   759 => x"c248ccf5",
   760 => x"cc78e6e5",
   761 => x"ccf5c087",
   762 => x"e0c048bf",
   763 => x"d0f5c080",
   764 => x"e2e5c258",
   765 => x"80c148bf",
   766 => x"58e6e5c2",
   767 => x"000d4c27",
   768 => x"bf97bf00",
   769 => x"c2029d4d",
   770 => x"e5c387e3",
   771 => x"dcc202ad",
   772 => x"ccf5c087",
   773 => x"a3cb4bbf",
   774 => x"cf4c1149",
   775 => x"d2c105ac",
   776 => x"df497587",
   777 => x"cd89c199",
   778 => x"f6edc291",
   779 => x"4aa3c181",
   780 => x"a3c35112",
   781 => x"c551124a",
   782 => x"51124aa3",
   783 => x"124aa3c7",
   784 => x"4aa3c951",
   785 => x"a3ce5112",
   786 => x"d051124a",
   787 => x"51124aa3",
   788 => x"124aa3d2",
   789 => x"4aa3d451",
   790 => x"a3d65112",
   791 => x"d851124a",
   792 => x"51124aa3",
   793 => x"124aa3dc",
   794 => x"4aa3de51",
   795 => x"7ec15112",
   796 => x"7487fac0",
   797 => x"0599c849",
   798 => x"7487ebc0",
   799 => x"0599d049",
   800 => x"66dc87d1",
   801 => x"87cbc002",
   802 => x"66dc4973",
   803 => x"0298700f",
   804 => x"6e87d3c0",
   805 => x"87c6c005",
   806 => x"48f6edc2",
   807 => x"f5c050c0",
   808 => x"c248bfcc",
   809 => x"eec287e1",
   810 => x"50c048c3",
   811 => x"f2edc27e",
   812 => x"e5c249bf",
   813 => x"714abfe2",
   814 => x"f6fb04aa",
   815 => x"d3f2c287",
   816 => x"c8c005bf",
   817 => x"eeedc287",
   818 => x"f8c102bf",
   819 => x"dee5c287",
   820 => x"fee849bf",
   821 => x"c2497087",
   822 => x"c459e2e5",
   823 => x"e5c248a6",
   824 => x"c278bfde",
   825 => x"02bfeeed",
   826 => x"c487d8c0",
   827 => x"ffcf4966",
   828 => x"99f8ffff",
   829 => x"c5c002a9",
   830 => x"c04cc087",
   831 => x"4cc187e1",
   832 => x"c487dcc0",
   833 => x"ffcf4966",
   834 => x"02a999f8",
   835 => x"c887c8c0",
   836 => x"78c048a6",
   837 => x"c887c5c0",
   838 => x"78c148a6",
   839 => x"744c66c8",
   840 => x"e0c0059c",
   841 => x"4966c487",
   842 => x"edc289c2",
   843 => x"914abfe6",
   844 => x"bffff1c2",
   845 => x"dae5c24a",
   846 => x"78a17248",
   847 => x"48e2e5c2",
   848 => x"def978c0",
   849 => x"f448c087",
   850 => x"87ffe68e",
   851 => x"00000000",
   852 => x"ffffffff",
   853 => x"00000d5c",
   854 => x"00000d65",
   855 => x"33544146",
   856 => x"20202032",
   857 => x"54414600",
   858 => x"20203631",
   859 => x"c21e0020",
   860 => x"48bfd8f2",
   861 => x"c905a8dd",
   862 => x"e1c2c187",
   863 => x"4a497087",
   864 => x"d4ff87c8",
   865 => x"78ffc348",
   866 => x"48724a68",
   867 => x"c21e4f26",
   868 => x"48bfd8f2",
   869 => x"c605a8dd",
   870 => x"edc1c187",
   871 => x"ff87d987",
   872 => x"ffc348d4",
   873 => x"48d0ff78",
   874 => x"ff78e1c0",
   875 => x"78d448d4",
   876 => x"48d7f2c2",
   877 => x"50bfd4ff",
   878 => x"ff1e4f26",
   879 => x"e0c048d0",
   880 => x"1e4f2678",
   881 => x"7087e7fe",
   882 => x"c6029949",
   883 => x"a9fbc087",
   884 => x"7187f105",
   885 => x"0e4f2648",
   886 => x"0e5c5b5e",
   887 => x"4cc04b71",
   888 => x"7087cbfe",
   889 => x"c0029949",
   890 => x"ecc087f9",
   891 => x"f2c002a9",
   892 => x"a9fbc087",
   893 => x"87ebc002",
   894 => x"acb766cc",
   895 => x"d087c703",
   896 => x"87c20266",
   897 => x"99715371",
   898 => x"c187c202",
   899 => x"87defd84",
   900 => x"02994970",
   901 => x"ecc087cd",
   902 => x"87c702a9",
   903 => x"05a9fbc0",
   904 => x"d087d5ff",
   905 => x"87c30266",
   906 => x"c07b97c0",
   907 => x"c405a9ec",
   908 => x"c54a7487",
   909 => x"c04a7487",
   910 => x"48728a0a",
   911 => x"4d2687c2",
   912 => x"4b264c26",
   913 => x"fc1e4f26",
   914 => x"497087e4",
   915 => x"aaf0c04a",
   916 => x"c087c904",
   917 => x"c301aaf9",
   918 => x"8af0c087",
   919 => x"04aac1c1",
   920 => x"dac187c9",
   921 => x"87c301aa",
   922 => x"728af7c0",
   923 => x"0e4f2648",
   924 => x"0e5c5b5e",
   925 => x"d4ff4a71",
   926 => x"c049724c",
   927 => x"4b7087e9",
   928 => x"87c2029b",
   929 => x"d0ff8bc1",
   930 => x"c178c548",
   931 => x"49737cd5",
   932 => x"e7c131c6",
   933 => x"4abf97d0",
   934 => x"70b07148",
   935 => x"48d0ff7c",
   936 => x"487378c4",
   937 => x"0e87d9fe",
   938 => x"5d5c5b5e",
   939 => x"7186f80e",
   940 => x"c07ec04b",
   941 => x"bf97cdfe",
   942 => x"c0059949",
   943 => x"a3c887ee",
   944 => x"49699749",
   945 => x"05a9c1c1",
   946 => x"a3c987dd",
   947 => x"49699749",
   948 => x"05a9d2c1",
   949 => x"a3ca87d1",
   950 => x"49699749",
   951 => x"05a9c3c1",
   952 => x"48df87c5",
   953 => x"c087e1c2",
   954 => x"87dcc248",
   955 => x"c087dffa",
   956 => x"cdfec04c",
   957 => x"c049bf97",
   958 => x"87cf04a9",
   959 => x"c187c4fb",
   960 => x"cdfec084",
   961 => x"ac49bf97",
   962 => x"c087f106",
   963 => x"bf97cdfe",
   964 => x"f987cf02",
   965 => x"497087d8",
   966 => x"87c60299",
   967 => x"05a9ecc0",
   968 => x"4cc087f1",
   969 => x"7087c7f9",
   970 => x"87c2f94d",
   971 => x"f858a6c8",
   972 => x"4a7087fc",
   973 => x"a3c884c1",
   974 => x"49699749",
   975 => x"87c702ad",
   976 => x"05adffc0",
   977 => x"c987e7c0",
   978 => x"699749a3",
   979 => x"a966c449",
   980 => x"4887c702",
   981 => x"05a8ffc0",
   982 => x"a3ca87d4",
   983 => x"49699749",
   984 => x"87c602aa",
   985 => x"05aaffc0",
   986 => x"7ec187c4",
   987 => x"ecc087d0",
   988 => x"87c602ad",
   989 => x"05adfbc0",
   990 => x"4cc087c4",
   991 => x"026e7ec1",
   992 => x"f887e1fe",
   993 => x"487487f4",
   994 => x"f1fa8ef8",
   995 => x"5e0e0087",
   996 => x"0e5d5c5b",
   997 => x"4d7186f8",
   998 => x"754bd4ff",
   999 => x"dcf2c21e",
  1000 => x"e0dfff49",
  1001 => x"7086c487",
  1002 => x"fbc40298",
  1003 => x"d2e7c187",
  1004 => x"49757ebf",
  1005 => x"de87f8fa",
  1006 => x"ebc005a8",
  1007 => x"c0497587",
  1008 => x"7087f9f6",
  1009 => x"87db0298",
  1010 => x"bfc0f7c2",
  1011 => x"49e1c01e",
  1012 => x"87c8f4c0",
  1013 => x"e7c186c4",
  1014 => x"50c048d0",
  1015 => x"49ccf7c2",
  1016 => x"c187ebfe",
  1017 => x"87c2c448",
  1018 => x"c548d0ff",
  1019 => x"7bd6c178",
  1020 => x"a2754ac0",
  1021 => x"c17b1149",
  1022 => x"aab7cb82",
  1023 => x"cc87f304",
  1024 => x"7bffc34a",
  1025 => x"e0c082c1",
  1026 => x"f404aab7",
  1027 => x"48d0ff87",
  1028 => x"ffc378c4",
  1029 => x"c178c57b",
  1030 => x"7bc17bd3",
  1031 => x"486e78c4",
  1032 => x"06a8b7c0",
  1033 => x"c287f0c2",
  1034 => x"4cbfe4f2",
  1035 => x"8874486e",
  1036 => x"9c747e70",
  1037 => x"87fdc102",
  1038 => x"4de6e5c2",
  1039 => x"c848a6c4",
  1040 => x"c08c78c0",
  1041 => x"c603acb7",
  1042 => x"a4c0c887",
  1043 => x"c24cc078",
  1044 => x"bf97d7f2",
  1045 => x"0299d049",
  1046 => x"1ec087d1",
  1047 => x"49dcf2c2",
  1048 => x"c487d5e1",
  1049 => x"4a497086",
  1050 => x"c287eec0",
  1051 => x"c21ee6e5",
  1052 => x"e149dcf2",
  1053 => x"86c487c2",
  1054 => x"ff4a4970",
  1055 => x"c5c848d0",
  1056 => x"7bd4c178",
  1057 => x"66c47b15",
  1058 => x"c888c148",
  1059 => x"987058a6",
  1060 => x"87f0ff05",
  1061 => x"c448d0ff",
  1062 => x"059a7278",
  1063 => x"48c087c5",
  1064 => x"c187c7c1",
  1065 => x"dcf2c21e",
  1066 => x"f1deff49",
  1067 => x"7486c487",
  1068 => x"c3fe059c",
  1069 => x"c0486e87",
  1070 => x"d106a8b7",
  1071 => x"dcf2c287",
  1072 => x"d078c048",
  1073 => x"f478c080",
  1074 => x"e8f2c280",
  1075 => x"486e78bf",
  1076 => x"01a8b7c0",
  1077 => x"ff87d0fd",
  1078 => x"78c548d0",
  1079 => x"c07bd3c1",
  1080 => x"c178c47b",
  1081 => x"87c2c048",
  1082 => x"8ef848c0",
  1083 => x"4c264d26",
  1084 => x"4f264b26",
  1085 => x"5c5b5e0e",
  1086 => x"711e0e5d",
  1087 => x"4d4cc04b",
  1088 => x"e8c004ab",
  1089 => x"e7fac087",
  1090 => x"029d751e",
  1091 => x"4ac087c4",
  1092 => x"4ac187c2",
  1093 => x"dbe94972",
  1094 => x"7086c487",
  1095 => x"6e84c17e",
  1096 => x"7387c205",
  1097 => x"7385c14c",
  1098 => x"d8ff06ac",
  1099 => x"26486e87",
  1100 => x"1e87f9fe",
  1101 => x"66c44a71",
  1102 => x"7287c505",
  1103 => x"87cef949",
  1104 => x"5e0e4f26",
  1105 => x"0e5d5c5b",
  1106 => x"494c711e",
  1107 => x"f3c291de",
  1108 => x"85714dc4",
  1109 => x"c1026d97",
  1110 => x"f2c287dc",
  1111 => x"744abff0",
  1112 => x"fe497282",
  1113 => x"7e7087ce",
  1114 => x"f2c0026e",
  1115 => x"f8f2c287",
  1116 => x"cb4a6e4b",
  1117 => x"effcfe49",
  1118 => x"cb4b7487",
  1119 => x"e4e7c193",
  1120 => x"c183c483",
  1121 => x"747bfac6",
  1122 => x"d0cbc149",
  1123 => x"c17b7587",
  1124 => x"bf97d1e7",
  1125 => x"f2c21e49",
  1126 => x"d6fe49f8",
  1127 => x"7486c487",
  1128 => x"f8cac149",
  1129 => x"c149c087",
  1130 => x"c287d7cc",
  1131 => x"c048d8f2",
  1132 => x"dd49c178",
  1133 => x"fc2687d9",
  1134 => x"6f4c87f2",
  1135 => x"6e696461",
  1136 => x"2e2e2e67",
  1137 => x"5b5e0e00",
  1138 => x"4b710e5c",
  1139 => x"f0f2c24a",
  1140 => x"497282bf",
  1141 => x"7087ddfc",
  1142 => x"c4029c4c",
  1143 => x"dbe54987",
  1144 => x"f0f2c287",
  1145 => x"c178c048",
  1146 => x"87e3dc49",
  1147 => x"0e87fffb",
  1148 => x"5d5c5b5e",
  1149 => x"c286f40e",
  1150 => x"c04de6e5",
  1151 => x"48a6c44c",
  1152 => x"f2c278c0",
  1153 => x"c049bff0",
  1154 => x"c1c106a9",
  1155 => x"e6e5c287",
  1156 => x"c0029848",
  1157 => x"fac087f8",
  1158 => x"66c81ee7",
  1159 => x"c487c702",
  1160 => x"78c048a6",
  1161 => x"a6c487c5",
  1162 => x"c478c148",
  1163 => x"c3e54966",
  1164 => x"7086c487",
  1165 => x"c484c14d",
  1166 => x"80c14866",
  1167 => x"c258a6c8",
  1168 => x"49bff0f2",
  1169 => x"87c603ac",
  1170 => x"ff059d75",
  1171 => x"4cc087c8",
  1172 => x"c3029d75",
  1173 => x"fac087e0",
  1174 => x"66c81ee7",
  1175 => x"cc87c702",
  1176 => x"78c048a6",
  1177 => x"a6cc87c5",
  1178 => x"cc78c148",
  1179 => x"c3e44966",
  1180 => x"7086c487",
  1181 => x"c2026e7e",
  1182 => x"496e87e9",
  1183 => x"699781cb",
  1184 => x"0299d049",
  1185 => x"c187d6c1",
  1186 => x"744ac5c7",
  1187 => x"c191cb49",
  1188 => x"7281e4e7",
  1189 => x"c381c879",
  1190 => x"497451ff",
  1191 => x"f3c291de",
  1192 => x"85714dc4",
  1193 => x"7d97c1c2",
  1194 => x"c049a5c1",
  1195 => x"edc251e0",
  1196 => x"02bf97f6",
  1197 => x"84c187d2",
  1198 => x"c24ba5c2",
  1199 => x"db4af6ed",
  1200 => x"e3f7fe49",
  1201 => x"87dbc187",
  1202 => x"c049a5cd",
  1203 => x"c284c151",
  1204 => x"4a6e4ba5",
  1205 => x"f7fe49cb",
  1206 => x"c6c187ce",
  1207 => x"c2c5c187",
  1208 => x"cb49744a",
  1209 => x"e4e7c191",
  1210 => x"c2797281",
  1211 => x"bf97f6ed",
  1212 => x"7487d802",
  1213 => x"c191de49",
  1214 => x"c4f3c284",
  1215 => x"c283714b",
  1216 => x"dd4af6ed",
  1217 => x"dff6fe49",
  1218 => x"7487d887",
  1219 => x"c293de4b",
  1220 => x"cb83c4f3",
  1221 => x"51c049a3",
  1222 => x"6e7384c1",
  1223 => x"fe49cb4a",
  1224 => x"c487c5f6",
  1225 => x"80c14866",
  1226 => x"c758a6c8",
  1227 => x"c5c003ac",
  1228 => x"fc056e87",
  1229 => x"487487e0",
  1230 => x"eff68ef4",
  1231 => x"1e731e87",
  1232 => x"cb494b71",
  1233 => x"e4e7c191",
  1234 => x"4aa1c881",
  1235 => x"48d0e7c1",
  1236 => x"a1c95012",
  1237 => x"cdfec04a",
  1238 => x"ca501248",
  1239 => x"d1e7c181",
  1240 => x"c1501148",
  1241 => x"bf97d1e7",
  1242 => x"49c01e49",
  1243 => x"c287c4f7",
  1244 => x"de48d8f2",
  1245 => x"d649c178",
  1246 => x"f52687d5",
  1247 => x"711e87f2",
  1248 => x"91cb494a",
  1249 => x"81e4e7c1",
  1250 => x"481181c8",
  1251 => x"58dcf2c2",
  1252 => x"48f0f2c2",
  1253 => x"49c178c0",
  1254 => x"2687f4d5",
  1255 => x"49c01e4f",
  1256 => x"87dec4c1",
  1257 => x"711e4f26",
  1258 => x"87d20299",
  1259 => x"48f9e8c1",
  1260 => x"80f750c0",
  1261 => x"40fecdc1",
  1262 => x"78dde7c1",
  1263 => x"e8c187ce",
  1264 => x"e7c148f5",
  1265 => x"80fc78d6",
  1266 => x"78ddcec1",
  1267 => x"5e0e4f26",
  1268 => x"710e5c5b",
  1269 => x"92cb4a4c",
  1270 => x"82e4e7c1",
  1271 => x"c949a2c8",
  1272 => x"6b974ba2",
  1273 => x"69971e4b",
  1274 => x"82ca1e49",
  1275 => x"e5c04912",
  1276 => x"49c087ca",
  1277 => x"7487d8d4",
  1278 => x"e0c1c149",
  1279 => x"f38ef887",
  1280 => x"731e87ec",
  1281 => x"494b711e",
  1282 => x"7387c3ff",
  1283 => x"87fefe49",
  1284 => x"1e87ddf3",
  1285 => x"4b711e73",
  1286 => x"024aa3c6",
  1287 => x"8ac187db",
  1288 => x"8a87d602",
  1289 => x"87dac102",
  1290 => x"fcc0028a",
  1291 => x"c0028a87",
  1292 => x"028a87e1",
  1293 => x"dbc187cb",
  1294 => x"fd49c787",
  1295 => x"dec187c0",
  1296 => x"f0f2c287",
  1297 => x"cbc102bf",
  1298 => x"88c14887",
  1299 => x"58f4f2c2",
  1300 => x"c287c1c1",
  1301 => x"02bff4f2",
  1302 => x"c287f9c0",
  1303 => x"48bff0f2",
  1304 => x"f2c280c1",
  1305 => x"ebc058f4",
  1306 => x"f0f2c287",
  1307 => x"89c649bf",
  1308 => x"59f4f2c2",
  1309 => x"03a9b7c0",
  1310 => x"f2c287da",
  1311 => x"78c048f0",
  1312 => x"f2c287d2",
  1313 => x"cb02bff4",
  1314 => x"f0f2c287",
  1315 => x"80c648bf",
  1316 => x"58f4f2c2",
  1317 => x"f6d149c0",
  1318 => x"c0497387",
  1319 => x"f187fefe",
  1320 => x"731e87ce",
  1321 => x"c24b711e",
  1322 => x"dd48d8f2",
  1323 => x"d149c078",
  1324 => x"497387dd",
  1325 => x"87e5fec0",
  1326 => x"0e87f5f0",
  1327 => x"5d5c5b5e",
  1328 => x"86ccff0e",
  1329 => x"c859a6d8",
  1330 => x"78c048a6",
  1331 => x"c8c180c4",
  1332 => x"80c47866",
  1333 => x"f2c278c1",
  1334 => x"78c148f4",
  1335 => x"bfd8f2c2",
  1336 => x"05a8de48",
  1337 => x"c6f487cb",
  1338 => x"cc497087",
  1339 => x"d0cf59a6",
  1340 => x"87dae287",
  1341 => x"e187cce3",
  1342 => x"4c7087f4",
  1343 => x"c10566d4",
  1344 => x"c4c187fc",
  1345 => x"80c44866",
  1346 => x"a6c47e70",
  1347 => x"78bf6e48",
  1348 => x"e3c11e72",
  1349 => x"66c848f6",
  1350 => x"4aa1c849",
  1351 => x"aa714120",
  1352 => x"1087f905",
  1353 => x"c14a2651",
  1354 => x"c14866c4",
  1355 => x"6e78fdcc",
  1356 => x"81c749bf",
  1357 => x"c4c15174",
  1358 => x"81c84966",
  1359 => x"c4c151c1",
  1360 => x"81c94966",
  1361 => x"c4c151c0",
  1362 => x"81ca4966",
  1363 => x"fbc051c0",
  1364 => x"87cf02ac",
  1365 => x"1ed81ec1",
  1366 => x"49bf66c8",
  1367 => x"f6e181c8",
  1368 => x"c186c887",
  1369 => x"c04866c8",
  1370 => x"87c701a8",
  1371 => x"c148a6c8",
  1372 => x"c187ce78",
  1373 => x"c14866c8",
  1374 => x"58a6d088",
  1375 => x"c2e187c3",
  1376 => x"48a6d887",
  1377 => x"9c7478c2",
  1378 => x"87f1cc02",
  1379 => x"c14866c8",
  1380 => x"03a866cc",
  1381 => x"dc87e6cc",
  1382 => x"78c048a6",
  1383 => x"78c080c4",
  1384 => x"87cadfff",
  1385 => x"66d44c70",
  1386 => x"05a8dd48",
  1387 => x"e0c087c7",
  1388 => x"66d448a6",
  1389 => x"acd0c178",
  1390 => x"87ebc005",
  1391 => x"87eedeff",
  1392 => x"87eadeff",
  1393 => x"ecc04c70",
  1394 => x"87c605ac",
  1395 => x"87f3dfff",
  1396 => x"d0c14c70",
  1397 => x"87c805ac",
  1398 => x"c14866d0",
  1399 => x"58a6d480",
  1400 => x"02acd0c1",
  1401 => x"c087d5ff",
  1402 => x"d448a6e4",
  1403 => x"e0c07866",
  1404 => x"e4c04866",
  1405 => x"ca05a866",
  1406 => x"e8c087d5",
  1407 => x"78c048a6",
  1408 => x"c080dcff",
  1409 => x"c04d7478",
  1410 => x"c9028dfb",
  1411 => x"8dc987db",
  1412 => x"c287db02",
  1413 => x"f7c1028d",
  1414 => x"028dc987",
  1415 => x"c487d8c4",
  1416 => x"c1c1028d",
  1417 => x"028dc187",
  1418 => x"c887ccc4",
  1419 => x"66c887f5",
  1420 => x"c191cb49",
  1421 => x"c48166c4",
  1422 => x"7e6a4aa1",
  1423 => x"e4c11e71",
  1424 => x"66c448c2",
  1425 => x"4aa1cc49",
  1426 => x"aa714120",
  1427 => x"87f8ff05",
  1428 => x"49265110",
  1429 => x"79e2d2c1",
  1430 => x"87d2dcff",
  1431 => x"a6c44c70",
  1432 => x"c878c148",
  1433 => x"a6dc87c3",
  1434 => x"78f0c048",
  1435 => x"87fedbff",
  1436 => x"ecc04c70",
  1437 => x"c4c002ac",
  1438 => x"a6e0c087",
  1439 => x"acecc05c",
  1440 => x"ff87cd02",
  1441 => x"7087e7db",
  1442 => x"acecc04c",
  1443 => x"87f3ff05",
  1444 => x"02acecc0",
  1445 => x"ff87c4c0",
  1446 => x"c087d3db",
  1447 => x"d01eca1e",
  1448 => x"91cb4966",
  1449 => x"4866ccc1",
  1450 => x"a6cc8071",
  1451 => x"4866c858",
  1452 => x"a6d080c4",
  1453 => x"bf66cc58",
  1454 => x"dadcff49",
  1455 => x"de1ec187",
  1456 => x"bf66d41e",
  1457 => x"cedcff49",
  1458 => x"7086d087",
  1459 => x"8909c049",
  1460 => x"59a6f0c0",
  1461 => x"4866ecc0",
  1462 => x"c006a8c0",
  1463 => x"ecc087ee",
  1464 => x"a8dd4866",
  1465 => x"87e4c003",
  1466 => x"49bf66c4",
  1467 => x"8166ecc0",
  1468 => x"c051e0c0",
  1469 => x"c14966ec",
  1470 => x"bf66c481",
  1471 => x"51c1c281",
  1472 => x"4966ecc0",
  1473 => x"66c481c2",
  1474 => x"51c081bf",
  1475 => x"ccc1486e",
  1476 => x"496e78fd",
  1477 => x"66d881c8",
  1478 => x"c9496e51",
  1479 => x"5166d081",
  1480 => x"81ca496e",
  1481 => x"d85166dc",
  1482 => x"80c14866",
  1483 => x"4858a6dc",
  1484 => x"78c180ec",
  1485 => x"ff87f2c4",
  1486 => x"7087cbdc",
  1487 => x"a6f0c049",
  1488 => x"c1dcff59",
  1489 => x"c0497087",
  1490 => x"dc59a6e0",
  1491 => x"ecc04866",
  1492 => x"cac005a8",
  1493 => x"48a6dc87",
  1494 => x"7866ecc0",
  1495 => x"ff87c4c0",
  1496 => x"c887cbd8",
  1497 => x"91cb4966",
  1498 => x"4866c4c1",
  1499 => x"7e708071",
  1500 => x"82c84a6e",
  1501 => x"81ca496e",
  1502 => x"5166ecc0",
  1503 => x"c14966dc",
  1504 => x"66ecc081",
  1505 => x"7148c189",
  1506 => x"c1497030",
  1507 => x"7a977189",
  1508 => x"bfe0f6c2",
  1509 => x"66ecc049",
  1510 => x"4a6a9729",
  1511 => x"c0987148",
  1512 => x"6e58a6f4",
  1513 => x"a681c449",
  1514 => x"c0786948",
  1515 => x"c04866e4",
  1516 => x"02a866e0",
  1517 => x"dc87c8c0",
  1518 => x"78c048a6",
  1519 => x"dc87c5c0",
  1520 => x"78c148a6",
  1521 => x"c01e66dc",
  1522 => x"66cc1ee0",
  1523 => x"c6d8ff49",
  1524 => x"7086c887",
  1525 => x"acb7c04c",
  1526 => x"87dbc106",
  1527 => x"744866c4",
  1528 => x"58a6c880",
  1529 => x"7449e0c0",
  1530 => x"4b66c489",
  1531 => x"4affe3c1",
  1532 => x"f3e2fe71",
  1533 => x"4866c487",
  1534 => x"a6c880c2",
  1535 => x"66e8c058",
  1536 => x"c080c148",
  1537 => x"c058a6ec",
  1538 => x"c14966f0",
  1539 => x"02a97081",
  1540 => x"c087c5c0",
  1541 => x"87c2c04d",
  1542 => x"1e754dc1",
  1543 => x"c049a4c2",
  1544 => x"887148e0",
  1545 => x"cc1e4970",
  1546 => x"d6ff4966",
  1547 => x"86c887e9",
  1548 => x"01a8b7c0",
  1549 => x"c087c6ff",
  1550 => x"c00266e8",
  1551 => x"496e87d1",
  1552 => x"e8c081c9",
  1553 => x"486e5166",
  1554 => x"78cecfc1",
  1555 => x"6e87ccc0",
  1556 => x"c281c949",
  1557 => x"c1486e51",
  1558 => x"c478c2d0",
  1559 => x"78c148a6",
  1560 => x"ff87c6c0",
  1561 => x"7087dcd5",
  1562 => x"0266c44c",
  1563 => x"c887f5c0",
  1564 => x"66cc4866",
  1565 => x"cbc004a8",
  1566 => x"4866c887",
  1567 => x"a6cc80c1",
  1568 => x"87e0c058",
  1569 => x"c14866cc",
  1570 => x"58a6d088",
  1571 => x"c187d5c0",
  1572 => x"c005acc6",
  1573 => x"66d887c8",
  1574 => x"dc80c148",
  1575 => x"d4ff58a6",
  1576 => x"4c7087e1",
  1577 => x"c14866d0",
  1578 => x"58a6d480",
  1579 => x"c0029c74",
  1580 => x"66c887cb",
  1581 => x"66ccc148",
  1582 => x"daf304a8",
  1583 => x"f9d3ff87",
  1584 => x"4866c887",
  1585 => x"c003a8c7",
  1586 => x"f2c287e5",
  1587 => x"78c048f4",
  1588 => x"cb4966c8",
  1589 => x"66c4c191",
  1590 => x"4aa1c481",
  1591 => x"52c04a6a",
  1592 => x"4866c879",
  1593 => x"a6cc80c1",
  1594 => x"04a8c758",
  1595 => x"ff87dbff",
  1596 => x"dfff8ecc",
  1597 => x"6f4c87f6",
  1598 => x"2a206461",
  1599 => x"3a00202e",
  1600 => x"49440020",
  1601 => x"77532050",
  1602 => x"68637469",
  1603 => x"1e007365",
  1604 => x"4b711e73",
  1605 => x"87c6029b",
  1606 => x"48f0f2c2",
  1607 => x"1ec778c0",
  1608 => x"bff0f2c2",
  1609 => x"e7c11e49",
  1610 => x"f2c21ee4",
  1611 => x"ee49bfd8",
  1612 => x"86cc87c9",
  1613 => x"bfd8f2c2",
  1614 => x"87eae949",
  1615 => x"c8029b73",
  1616 => x"e4e7c187",
  1617 => x"e6edc049",
  1618 => x"e3deff87",
  1619 => x"cdc71e87",
  1620 => x"fe49c187",
  1621 => x"e5fe87f9",
  1622 => x"987087dc",
  1623 => x"fe87cd02",
  1624 => x"7087f5ec",
  1625 => x"87c40298",
  1626 => x"87c24ac1",
  1627 => x"9a724ac0",
  1628 => x"c087ce05",
  1629 => x"e2e6c11e",
  1630 => x"d0f9c049",
  1631 => x"fe86c487",
  1632 => x"f3fbc087",
  1633 => x"c11ec087",
  1634 => x"c049ede6",
  1635 => x"c087fef8",
  1636 => x"f9fdc01e",
  1637 => x"c0497087",
  1638 => x"c287f2f8",
  1639 => x"8ef887ff",
  1640 => x"44534f26",
  1641 => x"69616620",
  1642 => x"2e64656c",
  1643 => x"6f6f4200",
  1644 => x"676e6974",
  1645 => x"002e2e2e",
  1646 => x"f0f2c21e",
  1647 => x"c278c048",
  1648 => x"c048d8f2",
  1649 => x"87c5fe78",
  1650 => x"87e1fdc0",
  1651 => x"4f2648c0",
  1652 => x"00010000",
  1653 => x"20800000",
  1654 => x"74697845",
  1655 => x"42208000",
  1656 => x"006b6361",
  1657 => x"0000137e",
  1658 => x"00002cc4",
  1659 => x"7e000000",
  1660 => x"e2000013",
  1661 => x"0000002c",
  1662 => x"137e0000",
  1663 => x"2d000000",
  1664 => x"00000000",
  1665 => x"00137e00",
  1666 => x"002d1e00",
  1667 => x"00000000",
  1668 => x"0000137e",
  1669 => x"00002d3c",
  1670 => x"7e000000",
  1671 => x"5a000013",
  1672 => x"0000002d",
  1673 => x"137e0000",
  1674 => x"2d780000",
  1675 => x"00000000",
  1676 => x"00137e00",
  1677 => x"00000000",
  1678 => x"00000000",
  1679 => x"00001413",
  1680 => x"00000000",
  1681 => x"1e000000",
  1682 => x"c048f0fe",
  1683 => x"7909cd78",
  1684 => x"1e4f2609",
  1685 => x"bff0fe1e",
  1686 => x"2626487e",
  1687 => x"f0fe1e4f",
  1688 => x"2678c148",
  1689 => x"f0fe1e4f",
  1690 => x"2678c048",
  1691 => x"4a711e4f",
  1692 => x"265252c0",
  1693 => x"5b5e0e4f",
  1694 => x"f40e5d5c",
  1695 => x"974d7186",
  1696 => x"a5c17e6d",
  1697 => x"486c974c",
  1698 => x"6e58a6c8",
  1699 => x"a866c448",
  1700 => x"ff87c505",
  1701 => x"87e6c048",
  1702 => x"c287caff",
  1703 => x"6c9749a5",
  1704 => x"4ba3714b",
  1705 => x"974b6b97",
  1706 => x"486e7e6c",
  1707 => x"a6c880c1",
  1708 => x"cc98c758",
  1709 => x"977058a6",
  1710 => x"87e1fe7c",
  1711 => x"8ef44873",
  1712 => x"4c264d26",
  1713 => x"4f264b26",
  1714 => x"5c5b5e0e",
  1715 => x"7186f40e",
  1716 => x"4a66d84c",
  1717 => x"c29affc3",
  1718 => x"6c974ba4",
  1719 => x"49a17349",
  1720 => x"6c975172",
  1721 => x"c1486e7e",
  1722 => x"58a6c880",
  1723 => x"a6cc98c7",
  1724 => x"f4547058",
  1725 => x"87caff8e",
  1726 => x"e8fd1e1e",
  1727 => x"4abfe087",
  1728 => x"c0e0c049",
  1729 => x"87cb0299",
  1730 => x"f6c21e72",
  1731 => x"f7fe49d6",
  1732 => x"fc86c487",
  1733 => x"7e7087fd",
  1734 => x"2687c2fd",
  1735 => x"c21e4f26",
  1736 => x"fd49d6f6",
  1737 => x"ebc187c7",
  1738 => x"dafc49f8",
  1739 => x"87c7c487",
  1740 => x"ff1e4f26",
  1741 => x"e1c848d0",
  1742 => x"48d4ff78",
  1743 => x"66c478c5",
  1744 => x"c387c302",
  1745 => x"66c878e0",
  1746 => x"ff87c602",
  1747 => x"f0c348d4",
  1748 => x"48d4ff78",
  1749 => x"d0ff7871",
  1750 => x"78e1c848",
  1751 => x"2678e0c0",
  1752 => x"5b5e0e4f",
  1753 => x"4c710e5c",
  1754 => x"49d6f6c2",
  1755 => x"7087c6fc",
  1756 => x"aab7c04a",
  1757 => x"87e2c204",
  1758 => x"05aaf0c3",
  1759 => x"f0c187c9",
  1760 => x"78c148e6",
  1761 => x"c387c3c2",
  1762 => x"c905aae0",
  1763 => x"eaf0c187",
  1764 => x"c178c148",
  1765 => x"f0c187f4",
  1766 => x"c602bfea",
  1767 => x"a2c0c287",
  1768 => x"7287c24b",
  1769 => x"059c744b",
  1770 => x"f0c187d1",
  1771 => x"c11ebfe6",
  1772 => x"1ebfeaf0",
  1773 => x"f9fd4972",
  1774 => x"c186c887",
  1775 => x"02bfe6f0",
  1776 => x"7387e0c0",
  1777 => x"29b7c449",
  1778 => x"c6f2c191",
  1779 => x"cf4a7381",
  1780 => x"c192c29a",
  1781 => x"70307248",
  1782 => x"72baff4a",
  1783 => x"70986948",
  1784 => x"7387db79",
  1785 => x"29b7c449",
  1786 => x"c6f2c191",
  1787 => x"cf4a7381",
  1788 => x"c392c29a",
  1789 => x"70307248",
  1790 => x"b069484a",
  1791 => x"f0c17970",
  1792 => x"78c048ea",
  1793 => x"48e6f0c1",
  1794 => x"f6c278c0",
  1795 => x"e4f949d6",
  1796 => x"c04a7087",
  1797 => x"fd03aab7",
  1798 => x"48c087de",
  1799 => x"4d2687c2",
  1800 => x"4b264c26",
  1801 => x"00004f26",
  1802 => x"00000000",
  1803 => x"711e0000",
  1804 => x"ecfc494a",
  1805 => x"1e4f2687",
  1806 => x"49724ac0",
  1807 => x"f2c191c4",
  1808 => x"79c081c6",
  1809 => x"b7d082c1",
  1810 => x"87ee04aa",
  1811 => x"5e0e4f26",
  1812 => x"0e5d5c5b",
  1813 => x"ccf84d71",
  1814 => x"c44a7587",
  1815 => x"c1922ab7",
  1816 => x"7582c6f2",
  1817 => x"c29ccf4c",
  1818 => x"4b496a94",
  1819 => x"9bc32b74",
  1820 => x"307448c2",
  1821 => x"bcff4c70",
  1822 => x"98714874",
  1823 => x"dcf77a70",
  1824 => x"fe487387",
  1825 => x"000087d8",
  1826 => x"00000000",
  1827 => x"00000000",
  1828 => x"00000000",
  1829 => x"00000000",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00000000",
  1834 => x"00000000",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"ff1e0000",
  1842 => x"e1c848d0",
  1843 => x"ff487178",
  1844 => x"c47808d4",
  1845 => x"d4ff4866",
  1846 => x"4f267808",
  1847 => x"c44a711e",
  1848 => x"721e4966",
  1849 => x"87deff49",
  1850 => x"c048d0ff",
  1851 => x"262678e0",
  1852 => x"1e731e4f",
  1853 => x"66c84b71",
  1854 => x"4a731e49",
  1855 => x"49a2e0c1",
  1856 => x"2687d9ff",
  1857 => x"4d2687c4",
  1858 => x"4b264c26",
  1859 => x"ff1e4f26",
  1860 => x"ffc34ad4",
  1861 => x"48d0ff7a",
  1862 => x"de78e1c0",
  1863 => x"e0f6c27a",
  1864 => x"48497abf",
  1865 => x"7a7028c8",
  1866 => x"28d04871",
  1867 => x"48717a70",
  1868 => x"7a7028d8",
  1869 => x"c048d0ff",
  1870 => x"4f2678e0",
  1871 => x"5c5b5e0e",
  1872 => x"4c710e5d",
  1873 => x"bfe0f6c2",
  1874 => x"2b744b4d",
  1875 => x"c19b66d0",
  1876 => x"ab66d483",
  1877 => x"c087c204",
  1878 => x"d04a744b",
  1879 => x"31724966",
  1880 => x"9975b9ff",
  1881 => x"30724873",
  1882 => x"71484a70",
  1883 => x"e4f6c2b0",
  1884 => x"87dafe58",
  1885 => x"4c264d26",
  1886 => x"4f264b26",
  1887 => x"5c5b5e0e",
  1888 => x"711e0e5d",
  1889 => x"e4f6c24c",
  1890 => x"c04ac04b",
  1891 => x"ccfe49f4",
  1892 => x"1e7487e6",
  1893 => x"49e4f6c2",
  1894 => x"87e9e7fe",
  1895 => x"497086c4",
  1896 => x"eac00299",
  1897 => x"a61ec487",
  1898 => x"f6c21e4d",
  1899 => x"effe49e4",
  1900 => x"86c887c0",
  1901 => x"d6029870",
  1902 => x"c14a7587",
  1903 => x"c449c5f8",
  1904 => x"e5cafe4b",
  1905 => x"02987087",
  1906 => x"48c087ca",
  1907 => x"c087edc0",
  1908 => x"87e8c048",
  1909 => x"c187f3c0",
  1910 => x"987087c4",
  1911 => x"c087c802",
  1912 => x"987087fc",
  1913 => x"c287f805",
  1914 => x"02bfc4f7",
  1915 => x"f6c287cc",
  1916 => x"f7c248e0",
  1917 => x"fc78bfc4",
  1918 => x"48c187d4",
  1919 => x"264d2626",
  1920 => x"264b264c",
  1921 => x"52415b4f",
  1922 => x"c01e0043",
  1923 => x"e4f6c21e",
  1924 => x"f2ebfe49",
  1925 => x"fcf6c287",
  1926 => x"2678c048",
  1927 => x"5e0e4f26",
  1928 => x"0e5d5c5b",
  1929 => x"7ec086f4",
  1930 => x"bffcf6c2",
  1931 => x"a8b7c348",
  1932 => x"c287d103",
  1933 => x"48bffcf6",
  1934 => x"f7c280c1",
  1935 => x"fbc058c0",
  1936 => x"87d9c648",
  1937 => x"49e4f6c2",
  1938 => x"87faf0fe",
  1939 => x"b7c04c70",
  1940 => x"87c403ac",
  1941 => x"87c5c648",
  1942 => x"bffcf6c2",
  1943 => x"028ac34a",
  1944 => x"8ac187d8",
  1945 => x"87c7c502",
  1946 => x"f2c2028a",
  1947 => x"c1028a87",
  1948 => x"028a87cf",
  1949 => x"c587dec3",
  1950 => x"4dc087d9",
  1951 => x"755ca6c8",
  1952 => x"c192c44a",
  1953 => x"c282fbff",
  1954 => x"754cf8f6",
  1955 => x"4b6c9784",
  1956 => x"a3c14b49",
  1957 => x"816a7c97",
  1958 => x"a6cc4811",
  1959 => x"4866c458",
  1960 => x"02a866c8",
  1961 => x"97c087c3",
  1962 => x"0566c87c",
  1963 => x"f6c287c7",
  1964 => x"a5c448fc",
  1965 => x"c485c178",
  1966 => x"ff04adb7",
  1967 => x"d2c487c1",
  1968 => x"c8f7c287",
  1969 => x"b7c848bf",
  1970 => x"87cb01a8",
  1971 => x"c602acca",
  1972 => x"05accd87",
  1973 => x"c287f3c0",
  1974 => x"4bbfc8f7",
  1975 => x"03abb7c8",
  1976 => x"f7c287d2",
  1977 => x"817349cc",
  1978 => x"c151e0c0",
  1979 => x"abb7c883",
  1980 => x"87eeff04",
  1981 => x"48d4f7c2",
  1982 => x"c150d2c1",
  1983 => x"cdc150cf",
  1984 => x"e450c050",
  1985 => x"c378c380",
  1986 => x"f7c287c9",
  1987 => x"4849bfc8",
  1988 => x"f7c280c1",
  1989 => x"c44858cc",
  1990 => x"517481a0",
  1991 => x"c087f4c2",
  1992 => x"04acb7f0",
  1993 => x"f9c087da",
  1994 => x"d301acb7",
  1995 => x"c0f7c287",
  1996 => x"91ca49bf",
  1997 => x"f0c04a74",
  1998 => x"c0f7c28a",
  1999 => x"78a17248",
  2000 => x"c002acca",
  2001 => x"accd87c6",
  2002 => x"87c7c205",
  2003 => x"48fcf6c2",
  2004 => x"fec178c3",
  2005 => x"b7f0c087",
  2006 => x"87db04ac",
  2007 => x"acb7f9c0",
  2008 => x"87d3c001",
  2009 => x"bfc4f7c2",
  2010 => x"7491d049",
  2011 => x"8af0c04a",
  2012 => x"48c4f7c2",
  2013 => x"c178a172",
  2014 => x"04acb7c1",
  2015 => x"c187dbc0",
  2016 => x"01acb7c6",
  2017 => x"c287d3c0",
  2018 => x"49bfc4f7",
  2019 => x"4a7491d0",
  2020 => x"c28af7c0",
  2021 => x"7248c4f7",
  2022 => x"acca78a1",
  2023 => x"87c6c002",
  2024 => x"c005accd",
  2025 => x"f6c287ed",
  2026 => x"78c348fc",
  2027 => x"c087e4c0",
  2028 => x"c005ace2",
  2029 => x"fbc087c6",
  2030 => x"87d7c07e",
  2031 => x"c002acca",
  2032 => x"accd87c6",
  2033 => x"87c9c005",
  2034 => x"48fcf6c2",
  2035 => x"c2c078c3",
  2036 => x"6e7e7487",
  2037 => x"87d0f902",
  2038 => x"ffc3486e",
  2039 => x"f88ef499",
  2040 => x"4f4387db",
  2041 => x"003d464e",
  2042 => x"00444f4d",
  2043 => x"454d414e",
  2044 => x"46454400",
  2045 => x"544c5541",
  2046 => x"e200303d",
  2047 => x"e800001f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
