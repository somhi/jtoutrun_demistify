
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"fc",x"f7",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"fc",x"f7",x"c2"),
    14 => (x"48",x"fc",x"e4",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e9",x"e5"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"81",x"48",x"73",x"1e"),
    47 => (x"72",x"05",x"a9",x"73"),
    48 => (x"26",x"87",x"f9",x"53"),
    49 => (x"4a",x"71",x"1e",x"4f"),
    50 => (x"48",x"49",x"66",x"c4"),
    51 => (x"a6",x"c8",x"88",x"c1"),
    52 => (x"02",x"99",x"71",x"58"),
    53 => (x"d4",x"ff",x"87",x"d6"),
    54 => (x"78",x"ff",x"c3",x"48"),
    55 => (x"66",x"c4",x"52",x"68"),
    56 => (x"88",x"c1",x"48",x"49"),
    57 => (x"71",x"58",x"a6",x"c8"),
    58 => (x"87",x"ea",x"05",x"99"),
    59 => (x"73",x"1e",x"4f",x"26"),
    60 => (x"4b",x"d4",x"ff",x"1e"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"7b",x"ff",x"c3",x"4a"),
    63 => (x"32",x"c8",x"49",x"6b"),
    64 => (x"ff",x"c3",x"b1",x"72"),
    65 => (x"c8",x"4a",x"6b",x"7b"),
    66 => (x"c3",x"b2",x"71",x"31"),
    67 => (x"49",x"6b",x"7b",x"ff"),
    68 => (x"b1",x"72",x"32",x"c8"),
    69 => (x"87",x"c4",x"48",x"71"),
    70 => (x"4c",x"26",x"4d",x"26"),
    71 => (x"4f",x"26",x"4b",x"26"),
    72 => (x"5c",x"5b",x"5e",x"0e"),
    73 => (x"4a",x"71",x"0e",x"5d"),
    74 => (x"72",x"4c",x"d4",x"ff"),
    75 => (x"99",x"ff",x"c3",x"49"),
    76 => (x"e4",x"c2",x"7c",x"71"),
    77 => (x"c8",x"05",x"bf",x"fc"),
    78 => (x"48",x"66",x"d0",x"87"),
    79 => (x"a6",x"d4",x"30",x"c9"),
    80 => (x"49",x"66",x"d0",x"58"),
    81 => (x"ff",x"c3",x"29",x"d8"),
    82 => (x"d0",x"7c",x"71",x"99"),
    83 => (x"29",x"d0",x"49",x"66"),
    84 => (x"71",x"99",x"ff",x"c3"),
    85 => (x"49",x"66",x"d0",x"7c"),
    86 => (x"ff",x"c3",x"29",x"c8"),
    87 => (x"d0",x"7c",x"71",x"99"),
    88 => (x"ff",x"c3",x"49",x"66"),
    89 => (x"72",x"7c",x"71",x"99"),
    90 => (x"c3",x"29",x"d0",x"49"),
    91 => (x"7c",x"71",x"99",x"ff"),
    92 => (x"f0",x"c9",x"4b",x"6c"),
    93 => (x"ff",x"c3",x"4d",x"ff"),
    94 => (x"87",x"d0",x"05",x"ab"),
    95 => (x"6c",x"7c",x"ff",x"c3"),
    96 => (x"02",x"8d",x"c1",x"4b"),
    97 => (x"ff",x"c3",x"87",x"c6"),
    98 => (x"87",x"f0",x"02",x"ab"),
    99 => (x"c7",x"fe",x"48",x"73"),
   100 => (x"49",x"c0",x"1e",x"87"),
   101 => (x"c3",x"48",x"d4",x"ff"),
   102 => (x"81",x"c1",x"78",x"ff"),
   103 => (x"a9",x"b7",x"c8",x"c3"),
   104 => (x"26",x"87",x"f1",x"04"),
   105 => (x"1e",x"73",x"1e",x"4f"),
   106 => (x"f8",x"c4",x"87",x"e7"),
   107 => (x"1e",x"c0",x"4b",x"df"),
   108 => (x"c1",x"f0",x"ff",x"c0"),
   109 => (x"e7",x"fd",x"49",x"f7"),
   110 => (x"c1",x"86",x"c4",x"87"),
   111 => (x"ea",x"c0",x"05",x"a8"),
   112 => (x"48",x"d4",x"ff",x"87"),
   113 => (x"c1",x"78",x"ff",x"c3"),
   114 => (x"c0",x"c0",x"c0",x"c0"),
   115 => (x"e1",x"c0",x"1e",x"c0"),
   116 => (x"49",x"e9",x"c1",x"f0"),
   117 => (x"c4",x"87",x"c9",x"fd"),
   118 => (x"05",x"98",x"70",x"86"),
   119 => (x"d4",x"ff",x"87",x"ca"),
   120 => (x"78",x"ff",x"c3",x"48"),
   121 => (x"87",x"cb",x"48",x"c1"),
   122 => (x"c1",x"87",x"e6",x"fe"),
   123 => (x"fd",x"fe",x"05",x"8b"),
   124 => (x"fc",x"48",x"c0",x"87"),
   125 => (x"73",x"1e",x"87",x"e6"),
   126 => (x"48",x"d4",x"ff",x"1e"),
   127 => (x"d3",x"78",x"ff",x"c3"),
   128 => (x"c0",x"1e",x"c0",x"4b"),
   129 => (x"c1",x"c1",x"f0",x"ff"),
   130 => (x"87",x"d4",x"fc",x"49"),
   131 => (x"98",x"70",x"86",x"c4"),
   132 => (x"ff",x"87",x"ca",x"05"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"cb",x"48",x"c1",x"78"),
   135 => (x"87",x"f1",x"fd",x"87"),
   136 => (x"ff",x"05",x"8b",x"c1"),
   137 => (x"48",x"c0",x"87",x"db"),
   138 => (x"0e",x"87",x"f1",x"fb"),
   139 => (x"0e",x"5c",x"5b",x"5e"),
   140 => (x"fd",x"4c",x"d4",x"ff"),
   141 => (x"ea",x"c6",x"87",x"db"),
   142 => (x"f0",x"e1",x"c0",x"1e"),
   143 => (x"fb",x"49",x"c8",x"c1"),
   144 => (x"86",x"c4",x"87",x"de"),
   145 => (x"c8",x"02",x"a8",x"c1"),
   146 => (x"87",x"ea",x"fe",x"87"),
   147 => (x"e2",x"c1",x"48",x"c0"),
   148 => (x"87",x"da",x"fa",x"87"),
   149 => (x"ff",x"cf",x"49",x"70"),
   150 => (x"ea",x"c6",x"99",x"ff"),
   151 => (x"87",x"c8",x"02",x"a9"),
   152 => (x"c0",x"87",x"d3",x"fe"),
   153 => (x"87",x"cb",x"c1",x"48"),
   154 => (x"c0",x"7c",x"ff",x"c3"),
   155 => (x"f4",x"fc",x"4b",x"f1"),
   156 => (x"02",x"98",x"70",x"87"),
   157 => (x"c0",x"87",x"eb",x"c0"),
   158 => (x"f0",x"ff",x"c0",x"1e"),
   159 => (x"fa",x"49",x"fa",x"c1"),
   160 => (x"86",x"c4",x"87",x"de"),
   161 => (x"d9",x"05",x"98",x"70"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"ff",x"c3",x"49",x"6c"),
   164 => (x"7c",x"7c",x"7c",x"7c"),
   165 => (x"02",x"99",x"c0",x"c1"),
   166 => (x"48",x"c1",x"87",x"c4"),
   167 => (x"48",x"c0",x"87",x"d5"),
   168 => (x"ab",x"c2",x"87",x"d1"),
   169 => (x"c0",x"87",x"c4",x"05"),
   170 => (x"c1",x"87",x"c8",x"48"),
   171 => (x"fd",x"fe",x"05",x"8b"),
   172 => (x"f9",x"48",x"c0",x"87"),
   173 => (x"73",x"1e",x"87",x"e4"),
   174 => (x"fc",x"e4",x"c2",x"1e"),
   175 => (x"c7",x"78",x"c1",x"48"),
   176 => (x"48",x"d0",x"ff",x"4b"),
   177 => (x"c8",x"fb",x"78",x"c2"),
   178 => (x"48",x"d0",x"ff",x"87"),
   179 => (x"1e",x"c0",x"78",x"c3"),
   180 => (x"c1",x"d0",x"e5",x"c0"),
   181 => (x"c7",x"f9",x"49",x"c0"),
   182 => (x"c1",x"86",x"c4",x"87"),
   183 => (x"87",x"c1",x"05",x"a8"),
   184 => (x"05",x"ab",x"c2",x"4b"),
   185 => (x"48",x"c0",x"87",x"c5"),
   186 => (x"c1",x"87",x"f9",x"c0"),
   187 => (x"d0",x"ff",x"05",x"8b"),
   188 => (x"87",x"f7",x"fc",x"87"),
   189 => (x"58",x"c0",x"e5",x"c2"),
   190 => (x"cd",x"05",x"98",x"70"),
   191 => (x"c0",x"1e",x"c1",x"87"),
   192 => (x"d0",x"c1",x"f0",x"ff"),
   193 => (x"87",x"d8",x"f8",x"49"),
   194 => (x"d4",x"ff",x"86",x"c4"),
   195 => (x"78",x"ff",x"c3",x"48"),
   196 => (x"c2",x"87",x"fc",x"c2"),
   197 => (x"ff",x"58",x"c4",x"e5"),
   198 => (x"78",x"c2",x"48",x"d0"),
   199 => (x"c3",x"48",x"d4",x"ff"),
   200 => (x"48",x"c1",x"78",x"ff"),
   201 => (x"0e",x"87",x"f5",x"f7"),
   202 => (x"5d",x"5c",x"5b",x"5e"),
   203 => (x"c0",x"4b",x"71",x"0e"),
   204 => (x"cd",x"ee",x"c5",x"4c"),
   205 => (x"d4",x"ff",x"4a",x"df"),
   206 => (x"78",x"ff",x"c3",x"48"),
   207 => (x"fe",x"c3",x"49",x"68"),
   208 => (x"fd",x"c0",x"05",x"a9"),
   209 => (x"73",x"4d",x"70",x"87"),
   210 => (x"87",x"cc",x"02",x"9b"),
   211 => (x"73",x"1e",x"66",x"d0"),
   212 => (x"87",x"f1",x"f5",x"49"),
   213 => (x"87",x"d6",x"86",x"c4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"ff",x"c3",x"78",x"d1"),
   216 => (x"48",x"66",x"d0",x"7d"),
   217 => (x"a6",x"d4",x"88",x"c1"),
   218 => (x"05",x"98",x"70",x"58"),
   219 => (x"d4",x"ff",x"87",x"f0"),
   220 => (x"78",x"ff",x"c3",x"48"),
   221 => (x"05",x"9b",x"73",x"78"),
   222 => (x"d0",x"ff",x"87",x"c5"),
   223 => (x"c1",x"78",x"d0",x"48"),
   224 => (x"8a",x"c1",x"4c",x"4a"),
   225 => (x"87",x"ee",x"fe",x"05"),
   226 => (x"cb",x"f6",x"48",x"74"),
   227 => (x"1e",x"73",x"1e",x"87"),
   228 => (x"4b",x"c0",x"4a",x"71"),
   229 => (x"c3",x"48",x"d4",x"ff"),
   230 => (x"d0",x"ff",x"78",x"ff"),
   231 => (x"78",x"c3",x"c4",x"48"),
   232 => (x"c3",x"48",x"d4",x"ff"),
   233 => (x"1e",x"72",x"78",x"ff"),
   234 => (x"c1",x"f0",x"ff",x"c0"),
   235 => (x"ef",x"f5",x"49",x"d1"),
   236 => (x"70",x"86",x"c4",x"87"),
   237 => (x"87",x"d2",x"05",x"98"),
   238 => (x"cc",x"1e",x"c0",x"c8"),
   239 => (x"e6",x"fd",x"49",x"66"),
   240 => (x"70",x"86",x"c4",x"87"),
   241 => (x"48",x"d0",x"ff",x"4b"),
   242 => (x"48",x"73",x"78",x"c2"),
   243 => (x"0e",x"87",x"cd",x"f5"),
   244 => (x"5d",x"5c",x"5b",x"5e"),
   245 => (x"c0",x"1e",x"c0",x"0e"),
   246 => (x"c9",x"c1",x"f0",x"ff"),
   247 => (x"87",x"c0",x"f5",x"49"),
   248 => (x"e5",x"c2",x"1e",x"d2"),
   249 => (x"fe",x"fc",x"49",x"c4"),
   250 => (x"c0",x"86",x"c8",x"87"),
   251 => (x"d2",x"84",x"c1",x"4c"),
   252 => (x"f8",x"04",x"ac",x"b7"),
   253 => (x"c4",x"e5",x"c2",x"87"),
   254 => (x"c3",x"49",x"bf",x"97"),
   255 => (x"c0",x"c1",x"99",x"c0"),
   256 => (x"e7",x"c0",x"05",x"a9"),
   257 => (x"cb",x"e5",x"c2",x"87"),
   258 => (x"d0",x"49",x"bf",x"97"),
   259 => (x"cc",x"e5",x"c2",x"31"),
   260 => (x"c8",x"4a",x"bf",x"97"),
   261 => (x"c2",x"b1",x"72",x"32"),
   262 => (x"bf",x"97",x"cd",x"e5"),
   263 => (x"4c",x"71",x"b1",x"4a"),
   264 => (x"ff",x"ff",x"ff",x"cf"),
   265 => (x"ca",x"84",x"c1",x"9c"),
   266 => (x"87",x"e7",x"c1",x"34"),
   267 => (x"97",x"cd",x"e5",x"c2"),
   268 => (x"31",x"c1",x"49",x"bf"),
   269 => (x"e5",x"c2",x"99",x"c6"),
   270 => (x"4a",x"bf",x"97",x"ce"),
   271 => (x"72",x"2a",x"b7",x"c7"),
   272 => (x"c9",x"e5",x"c2",x"b1"),
   273 => (x"4d",x"4a",x"bf",x"97"),
   274 => (x"e5",x"c2",x"9d",x"cf"),
   275 => (x"4a",x"bf",x"97",x"ca"),
   276 => (x"32",x"ca",x"9a",x"c3"),
   277 => (x"97",x"cb",x"e5",x"c2"),
   278 => (x"33",x"c2",x"4b",x"bf"),
   279 => (x"e5",x"c2",x"b2",x"73"),
   280 => (x"4b",x"bf",x"97",x"cc"),
   281 => (x"c6",x"9b",x"c0",x"c3"),
   282 => (x"b2",x"73",x"2b",x"b7"),
   283 => (x"48",x"c1",x"81",x"c2"),
   284 => (x"49",x"70",x"30",x"71"),
   285 => (x"30",x"75",x"48",x"c1"),
   286 => (x"4c",x"72",x"4d",x"70"),
   287 => (x"94",x"71",x"84",x"c1"),
   288 => (x"ad",x"b7",x"c0",x"c8"),
   289 => (x"c1",x"87",x"cc",x"06"),
   290 => (x"c8",x"2d",x"b7",x"34"),
   291 => (x"01",x"ad",x"b7",x"c0"),
   292 => (x"74",x"87",x"f4",x"ff"),
   293 => (x"87",x"c0",x"f2",x"48"),
   294 => (x"5c",x"5b",x"5e",x"0e"),
   295 => (x"86",x"f8",x"0e",x"5d"),
   296 => (x"48",x"ea",x"ed",x"c2"),
   297 => (x"e5",x"c2",x"78",x"c0"),
   298 => (x"49",x"c0",x"1e",x"e2"),
   299 => (x"c4",x"87",x"de",x"fb"),
   300 => (x"05",x"98",x"70",x"86"),
   301 => (x"48",x"c0",x"87",x"c5"),
   302 => (x"c0",x"87",x"ce",x"c9"),
   303 => (x"c0",x"7e",x"c1",x"4d"),
   304 => (x"49",x"bf",x"d8",x"f5"),
   305 => (x"4a",x"d8",x"e6",x"c2"),
   306 => (x"ee",x"4b",x"c8",x"71"),
   307 => (x"98",x"70",x"87",x"dc"),
   308 => (x"c0",x"87",x"c2",x"05"),
   309 => (x"d4",x"f5",x"c0",x"7e"),
   310 => (x"e6",x"c2",x"49",x"bf"),
   311 => (x"c8",x"71",x"4a",x"f4"),
   312 => (x"87",x"c6",x"ee",x"4b"),
   313 => (x"c2",x"05",x"98",x"70"),
   314 => (x"6e",x"7e",x"c0",x"87"),
   315 => (x"87",x"fd",x"c0",x"02"),
   316 => (x"bf",x"e8",x"ec",x"c2"),
   317 => (x"e0",x"ed",x"c2",x"4d"),
   318 => (x"48",x"7e",x"bf",x"9f"),
   319 => (x"a8",x"ea",x"d6",x"c5"),
   320 => (x"c2",x"87",x"c7",x"05"),
   321 => (x"4d",x"bf",x"e8",x"ec"),
   322 => (x"48",x"6e",x"87",x"ce"),
   323 => (x"a8",x"d5",x"e9",x"ca"),
   324 => (x"c0",x"87",x"c5",x"02"),
   325 => (x"87",x"f1",x"c7",x"48"),
   326 => (x"1e",x"e2",x"e5",x"c2"),
   327 => (x"ec",x"f9",x"49",x"75"),
   328 => (x"70",x"86",x"c4",x"87"),
   329 => (x"87",x"c5",x"05",x"98"),
   330 => (x"dc",x"c7",x"48",x"c0"),
   331 => (x"d4",x"f5",x"c0",x"87"),
   332 => (x"e6",x"c2",x"49",x"bf"),
   333 => (x"c8",x"71",x"4a",x"f4"),
   334 => (x"87",x"ee",x"ec",x"4b"),
   335 => (x"c8",x"05",x"98",x"70"),
   336 => (x"ea",x"ed",x"c2",x"87"),
   337 => (x"da",x"78",x"c1",x"48"),
   338 => (x"d8",x"f5",x"c0",x"87"),
   339 => (x"e6",x"c2",x"49",x"bf"),
   340 => (x"c8",x"71",x"4a",x"d8"),
   341 => (x"87",x"d2",x"ec",x"4b"),
   342 => (x"c0",x"02",x"98",x"70"),
   343 => (x"48",x"c0",x"87",x"c5"),
   344 => (x"c2",x"87",x"e6",x"c6"),
   345 => (x"bf",x"97",x"e0",x"ed"),
   346 => (x"a9",x"d5",x"c1",x"49"),
   347 => (x"87",x"cd",x"c0",x"05"),
   348 => (x"97",x"e1",x"ed",x"c2"),
   349 => (x"ea",x"c2",x"49",x"bf"),
   350 => (x"c5",x"c0",x"02",x"a9"),
   351 => (x"c6",x"48",x"c0",x"87"),
   352 => (x"e5",x"c2",x"87",x"c7"),
   353 => (x"7e",x"bf",x"97",x"e2"),
   354 => (x"a8",x"e9",x"c3",x"48"),
   355 => (x"87",x"ce",x"c0",x"02"),
   356 => (x"eb",x"c3",x"48",x"6e"),
   357 => (x"c5",x"c0",x"02",x"a8"),
   358 => (x"c5",x"48",x"c0",x"87"),
   359 => (x"e5",x"c2",x"87",x"eb"),
   360 => (x"49",x"bf",x"97",x"ed"),
   361 => (x"cc",x"c0",x"05",x"99"),
   362 => (x"ee",x"e5",x"c2",x"87"),
   363 => (x"c2",x"49",x"bf",x"97"),
   364 => (x"c5",x"c0",x"02",x"a9"),
   365 => (x"c5",x"48",x"c0",x"87"),
   366 => (x"e5",x"c2",x"87",x"cf"),
   367 => (x"48",x"bf",x"97",x"ef"),
   368 => (x"58",x"e6",x"ed",x"c2"),
   369 => (x"c1",x"48",x"4c",x"70"),
   370 => (x"ea",x"ed",x"c2",x"88"),
   371 => (x"f0",x"e5",x"c2",x"58"),
   372 => (x"75",x"49",x"bf",x"97"),
   373 => (x"f1",x"e5",x"c2",x"81"),
   374 => (x"c8",x"4a",x"bf",x"97"),
   375 => (x"7e",x"a1",x"72",x"32"),
   376 => (x"48",x"f7",x"f1",x"c2"),
   377 => (x"e5",x"c2",x"78",x"6e"),
   378 => (x"48",x"bf",x"97",x"f2"),
   379 => (x"c2",x"58",x"a6",x"c8"),
   380 => (x"02",x"bf",x"ea",x"ed"),
   381 => (x"c0",x"87",x"d4",x"c2"),
   382 => (x"49",x"bf",x"d4",x"f5"),
   383 => (x"4a",x"f4",x"e6",x"c2"),
   384 => (x"e9",x"4b",x"c8",x"71"),
   385 => (x"98",x"70",x"87",x"e4"),
   386 => (x"87",x"c5",x"c0",x"02"),
   387 => (x"f8",x"c3",x"48",x"c0"),
   388 => (x"e2",x"ed",x"c2",x"87"),
   389 => (x"f2",x"c2",x"4c",x"bf"),
   390 => (x"e6",x"c2",x"5c",x"cb"),
   391 => (x"49",x"bf",x"97",x"c7"),
   392 => (x"e6",x"c2",x"31",x"c8"),
   393 => (x"4a",x"bf",x"97",x"c6"),
   394 => (x"e6",x"c2",x"49",x"a1"),
   395 => (x"4a",x"bf",x"97",x"c8"),
   396 => (x"a1",x"72",x"32",x"d0"),
   397 => (x"c9",x"e6",x"c2",x"49"),
   398 => (x"d8",x"4a",x"bf",x"97"),
   399 => (x"49",x"a1",x"72",x"32"),
   400 => (x"c2",x"91",x"66",x"c4"),
   401 => (x"81",x"bf",x"f7",x"f1"),
   402 => (x"59",x"ff",x"f1",x"c2"),
   403 => (x"97",x"cf",x"e6",x"c2"),
   404 => (x"32",x"c8",x"4a",x"bf"),
   405 => (x"97",x"ce",x"e6",x"c2"),
   406 => (x"4a",x"a2",x"4b",x"bf"),
   407 => (x"97",x"d0",x"e6",x"c2"),
   408 => (x"33",x"d0",x"4b",x"bf"),
   409 => (x"c2",x"4a",x"a2",x"73"),
   410 => (x"bf",x"97",x"d1",x"e6"),
   411 => (x"d8",x"9b",x"cf",x"4b"),
   412 => (x"4a",x"a2",x"73",x"33"),
   413 => (x"5a",x"c3",x"f2",x"c2"),
   414 => (x"bf",x"ff",x"f1",x"c2"),
   415 => (x"74",x"8a",x"c2",x"4a"),
   416 => (x"c3",x"f2",x"c2",x"92"),
   417 => (x"78",x"a1",x"72",x"48"),
   418 => (x"c2",x"87",x"ca",x"c1"),
   419 => (x"bf",x"97",x"f4",x"e5"),
   420 => (x"c2",x"31",x"c8",x"49"),
   421 => (x"bf",x"97",x"f3",x"e5"),
   422 => (x"c2",x"49",x"a1",x"4a"),
   423 => (x"c2",x"59",x"f2",x"ed"),
   424 => (x"49",x"bf",x"ee",x"ed"),
   425 => (x"ff",x"c7",x"31",x"c5"),
   426 => (x"c2",x"29",x"c9",x"81"),
   427 => (x"c2",x"59",x"cb",x"f2"),
   428 => (x"bf",x"97",x"f9",x"e5"),
   429 => (x"c2",x"32",x"c8",x"4a"),
   430 => (x"bf",x"97",x"f8",x"e5"),
   431 => (x"c4",x"4a",x"a2",x"4b"),
   432 => (x"82",x"6e",x"92",x"66"),
   433 => (x"5a",x"c7",x"f2",x"c2"),
   434 => (x"48",x"ff",x"f1",x"c2"),
   435 => (x"f1",x"c2",x"78",x"c0"),
   436 => (x"a1",x"72",x"48",x"fb"),
   437 => (x"cb",x"f2",x"c2",x"78"),
   438 => (x"ff",x"f1",x"c2",x"48"),
   439 => (x"f2",x"c2",x"78",x"bf"),
   440 => (x"f2",x"c2",x"48",x"cf"),
   441 => (x"c2",x"78",x"bf",x"c3"),
   442 => (x"02",x"bf",x"ea",x"ed"),
   443 => (x"74",x"87",x"c9",x"c0"),
   444 => (x"70",x"30",x"c4",x"48"),
   445 => (x"87",x"c9",x"c0",x"7e"),
   446 => (x"bf",x"c7",x"f2",x"c2"),
   447 => (x"70",x"30",x"c4",x"48"),
   448 => (x"ee",x"ed",x"c2",x"7e"),
   449 => (x"c1",x"78",x"6e",x"48"),
   450 => (x"26",x"8e",x"f8",x"48"),
   451 => (x"26",x"4c",x"26",x"4d"),
   452 => (x"0e",x"4f",x"26",x"4b"),
   453 => (x"5d",x"5c",x"5b",x"5e"),
   454 => (x"c2",x"4a",x"71",x"0e"),
   455 => (x"02",x"bf",x"ea",x"ed"),
   456 => (x"4b",x"72",x"87",x"cb"),
   457 => (x"4c",x"72",x"2b",x"c7"),
   458 => (x"c9",x"9c",x"ff",x"c1"),
   459 => (x"c8",x"4b",x"72",x"87"),
   460 => (x"c3",x"4c",x"72",x"2b"),
   461 => (x"f1",x"c2",x"9c",x"ff"),
   462 => (x"c0",x"83",x"bf",x"f7"),
   463 => (x"ab",x"bf",x"d0",x"f5"),
   464 => (x"c0",x"87",x"d9",x"02"),
   465 => (x"c2",x"5b",x"d4",x"f5"),
   466 => (x"73",x"1e",x"e2",x"e5"),
   467 => (x"87",x"fd",x"f0",x"49"),
   468 => (x"98",x"70",x"86",x"c4"),
   469 => (x"c0",x"87",x"c5",x"05"),
   470 => (x"87",x"e6",x"c0",x"48"),
   471 => (x"bf",x"ea",x"ed",x"c2"),
   472 => (x"74",x"87",x"d2",x"02"),
   473 => (x"c2",x"91",x"c4",x"49"),
   474 => (x"69",x"81",x"e2",x"e5"),
   475 => (x"ff",x"ff",x"cf",x"4d"),
   476 => (x"cb",x"9d",x"ff",x"ff"),
   477 => (x"c2",x"49",x"74",x"87"),
   478 => (x"e2",x"e5",x"c2",x"91"),
   479 => (x"4d",x"69",x"9f",x"81"),
   480 => (x"c6",x"fe",x"48",x"75"),
   481 => (x"5b",x"5e",x"0e",x"87"),
   482 => (x"f8",x"0e",x"5d",x"5c"),
   483 => (x"9c",x"4c",x"71",x"86"),
   484 => (x"c0",x"87",x"c5",x"05"),
   485 => (x"87",x"c1",x"c3",x"48"),
   486 => (x"6e",x"7e",x"a4",x"c8"),
   487 => (x"d8",x"78",x"c0",x"48"),
   488 => (x"87",x"c7",x"02",x"66"),
   489 => (x"bf",x"97",x"66",x"d8"),
   490 => (x"c0",x"87",x"c5",x"05"),
   491 => (x"87",x"e9",x"c2",x"48"),
   492 => (x"49",x"c1",x"1e",x"c0"),
   493 => (x"c4",x"87",x"fd",x"ce"),
   494 => (x"9d",x"4d",x"70",x"86"),
   495 => (x"87",x"c2",x"c1",x"02"),
   496 => (x"4a",x"f2",x"ed",x"c2"),
   497 => (x"e2",x"49",x"66",x"d8"),
   498 => (x"98",x"70",x"87",x"c5"),
   499 => (x"87",x"f2",x"c0",x"02"),
   500 => (x"66",x"d8",x"4a",x"75"),
   501 => (x"e2",x"4b",x"cb",x"49"),
   502 => (x"98",x"70",x"87",x"ea"),
   503 => (x"87",x"e2",x"c0",x"02"),
   504 => (x"9d",x"75",x"1e",x"c0"),
   505 => (x"c8",x"87",x"c7",x"02"),
   506 => (x"78",x"c0",x"48",x"a6"),
   507 => (x"a6",x"c8",x"87",x"c5"),
   508 => (x"c8",x"78",x"c1",x"48"),
   509 => (x"fb",x"cd",x"49",x"66"),
   510 => (x"70",x"86",x"c4",x"87"),
   511 => (x"fe",x"05",x"9d",x"4d"),
   512 => (x"9d",x"75",x"87",x"fe"),
   513 => (x"87",x"cf",x"c1",x"02"),
   514 => (x"6e",x"49",x"a5",x"dc"),
   515 => (x"da",x"78",x"69",x"48"),
   516 => (x"a6",x"c4",x"49",x"a5"),
   517 => (x"78",x"a4",x"c4",x"48"),
   518 => (x"c4",x"48",x"69",x"9f"),
   519 => (x"c2",x"78",x"08",x"66"),
   520 => (x"02",x"bf",x"ea",x"ed"),
   521 => (x"a5",x"d4",x"87",x"d2"),
   522 => (x"49",x"69",x"9f",x"49"),
   523 => (x"99",x"ff",x"ff",x"c0"),
   524 => (x"30",x"d0",x"48",x"71"),
   525 => (x"87",x"c2",x"7e",x"70"),
   526 => (x"49",x"6e",x"7e",x"c0"),
   527 => (x"bf",x"66",x"c4",x"48"),
   528 => (x"08",x"66",x"c4",x"80"),
   529 => (x"cc",x"7c",x"c0",x"78"),
   530 => (x"66",x"c4",x"49",x"a4"),
   531 => (x"a4",x"d0",x"79",x"bf"),
   532 => (x"c1",x"79",x"c0",x"49"),
   533 => (x"c0",x"87",x"c2",x"48"),
   534 => (x"fa",x"8e",x"f8",x"48"),
   535 => (x"5e",x"0e",x"87",x"ed"),
   536 => (x"0e",x"5d",x"5c",x"5b"),
   537 => (x"02",x"9c",x"4c",x"71"),
   538 => (x"c8",x"87",x"ca",x"c1"),
   539 => (x"02",x"69",x"49",x"a4"),
   540 => (x"d0",x"87",x"c2",x"c1"),
   541 => (x"49",x"6c",x"4a",x"66"),
   542 => (x"5a",x"a6",x"d4",x"82"),
   543 => (x"b9",x"4d",x"66",x"d0"),
   544 => (x"bf",x"e6",x"ed",x"c2"),
   545 => (x"72",x"ba",x"ff",x"4a"),
   546 => (x"02",x"99",x"71",x"99"),
   547 => (x"c4",x"87",x"e4",x"c0"),
   548 => (x"49",x"6b",x"4b",x"a4"),
   549 => (x"70",x"87",x"fc",x"f9"),
   550 => (x"e2",x"ed",x"c2",x"7b"),
   551 => (x"81",x"6c",x"49",x"bf"),
   552 => (x"b9",x"75",x"7c",x"71"),
   553 => (x"bf",x"e6",x"ed",x"c2"),
   554 => (x"72",x"ba",x"ff",x"4a"),
   555 => (x"05",x"99",x"71",x"99"),
   556 => (x"75",x"87",x"dc",x"ff"),
   557 => (x"87",x"d3",x"f9",x"7c"),
   558 => (x"71",x"1e",x"73",x"1e"),
   559 => (x"c7",x"02",x"9b",x"4b"),
   560 => (x"49",x"a3",x"c8",x"87"),
   561 => (x"87",x"c5",x"05",x"69"),
   562 => (x"f7",x"c0",x"48",x"c0"),
   563 => (x"fb",x"f1",x"c2",x"87"),
   564 => (x"a3",x"c4",x"4a",x"bf"),
   565 => (x"c2",x"49",x"69",x"49"),
   566 => (x"e2",x"ed",x"c2",x"89"),
   567 => (x"a2",x"71",x"91",x"bf"),
   568 => (x"e6",x"ed",x"c2",x"4a"),
   569 => (x"99",x"6b",x"49",x"bf"),
   570 => (x"c0",x"4a",x"a2",x"71"),
   571 => (x"c8",x"5a",x"d4",x"f5"),
   572 => (x"49",x"72",x"1e",x"66"),
   573 => (x"c4",x"87",x"d6",x"ea"),
   574 => (x"05",x"98",x"70",x"86"),
   575 => (x"48",x"c0",x"87",x"c4"),
   576 => (x"48",x"c1",x"87",x"c2"),
   577 => (x"0e",x"87",x"c8",x"f8"),
   578 => (x"0e",x"5c",x"5b",x"5e"),
   579 => (x"d0",x"4b",x"71",x"1e"),
   580 => (x"2c",x"c9",x"4c",x"66"),
   581 => (x"c1",x"02",x"9b",x"73"),
   582 => (x"a3",x"c8",x"87",x"d4"),
   583 => (x"c1",x"02",x"69",x"49"),
   584 => (x"ed",x"c2",x"87",x"cc"),
   585 => (x"ff",x"49",x"bf",x"e6"),
   586 => (x"99",x"4a",x"6b",x"b9"),
   587 => (x"03",x"ac",x"71",x"7e"),
   588 => (x"7b",x"c0",x"87",x"d1"),
   589 => (x"c0",x"49",x"a3",x"d0"),
   590 => (x"4a",x"a3",x"cc",x"79"),
   591 => (x"6a",x"49",x"a3",x"c4"),
   592 => (x"72",x"87",x"c2",x"79"),
   593 => (x"02",x"9c",x"74",x"8c"),
   594 => (x"49",x"87",x"e3",x"c0"),
   595 => (x"fc",x"49",x"73",x"1e"),
   596 => (x"86",x"c4",x"87",x"cc"),
   597 => (x"c7",x"49",x"66",x"d0"),
   598 => (x"cb",x"02",x"99",x"ff"),
   599 => (x"e2",x"e5",x"c2",x"87"),
   600 => (x"fd",x"49",x"73",x"1e"),
   601 => (x"86",x"c4",x"87",x"d2"),
   602 => (x"d0",x"49",x"a3",x"d0"),
   603 => (x"f6",x"26",x"79",x"66"),
   604 => (x"5e",x"0e",x"87",x"db"),
   605 => (x"0e",x"5d",x"5c",x"5b"),
   606 => (x"a6",x"d0",x"86",x"f0"),
   607 => (x"66",x"e4",x"c0",x"59"),
   608 => (x"02",x"66",x"cc",x"4b"),
   609 => (x"c8",x"48",x"87",x"ca"),
   610 => (x"6e",x"7e",x"70",x"80"),
   611 => (x"87",x"c5",x"05",x"bf"),
   612 => (x"ec",x"c3",x"48",x"c0"),
   613 => (x"4c",x"66",x"cc",x"87"),
   614 => (x"49",x"73",x"84",x"d0"),
   615 => (x"6c",x"48",x"a6",x"c4"),
   616 => (x"81",x"66",x"c4",x"78"),
   617 => (x"bf",x"6e",x"80",x"c4"),
   618 => (x"a9",x"66",x"c8",x"78"),
   619 => (x"49",x"87",x"c6",x"06"),
   620 => (x"71",x"89",x"66",x"c4"),
   621 => (x"ab",x"b7",x"c0",x"4b"),
   622 => (x"48",x"87",x"c4",x"01"),
   623 => (x"c4",x"87",x"c2",x"c3"),
   624 => (x"ff",x"c7",x"48",x"66"),
   625 => (x"6e",x"7e",x"70",x"98"),
   626 => (x"87",x"c9",x"c1",x"02"),
   627 => (x"6e",x"49",x"c0",x"c8"),
   628 => (x"c2",x"4a",x"71",x"89"),
   629 => (x"6e",x"4d",x"e2",x"e5"),
   630 => (x"aa",x"b7",x"73",x"85"),
   631 => (x"4a",x"87",x"c1",x"06"),
   632 => (x"c4",x"48",x"49",x"72"),
   633 => (x"7c",x"70",x"80",x"66"),
   634 => (x"c1",x"49",x"8b",x"72"),
   635 => (x"02",x"99",x"71",x"8a"),
   636 => (x"e0",x"c0",x"87",x"d9"),
   637 => (x"50",x"15",x"48",x"66"),
   638 => (x"48",x"66",x"e0",x"c0"),
   639 => (x"e4",x"c0",x"80",x"c1"),
   640 => (x"49",x"72",x"58",x"a6"),
   641 => (x"99",x"71",x"8a",x"c1"),
   642 => (x"c1",x"87",x"e7",x"05"),
   643 => (x"49",x"66",x"d0",x"1e"),
   644 => (x"c4",x"87",x"cb",x"f9"),
   645 => (x"ab",x"b7",x"c0",x"86"),
   646 => (x"87",x"e3",x"c1",x"06"),
   647 => (x"4d",x"66",x"e0",x"c0"),
   648 => (x"ab",x"b7",x"ff",x"c7"),
   649 => (x"87",x"e2",x"c0",x"06"),
   650 => (x"66",x"d0",x"1e",x"75"),
   651 => (x"87",x"c8",x"fa",x"49"),
   652 => (x"6c",x"85",x"c0",x"c8"),
   653 => (x"80",x"c0",x"c8",x"48"),
   654 => (x"c0",x"c8",x"7c",x"70"),
   655 => (x"d4",x"1e",x"c1",x"8b"),
   656 => (x"d9",x"f8",x"49",x"66"),
   657 => (x"c0",x"86",x"c8",x"87"),
   658 => (x"e5",x"c2",x"87",x"ee"),
   659 => (x"66",x"d0",x"1e",x"e2"),
   660 => (x"87",x"e4",x"f9",x"49"),
   661 => (x"e5",x"c2",x"86",x"c4"),
   662 => (x"49",x"73",x"4a",x"e2"),
   663 => (x"70",x"80",x"6c",x"48"),
   664 => (x"c1",x"49",x"73",x"7c"),
   665 => (x"02",x"99",x"71",x"8b"),
   666 => (x"97",x"12",x"87",x"ce"),
   667 => (x"73",x"85",x"c1",x"7d"),
   668 => (x"71",x"8b",x"c1",x"49"),
   669 => (x"87",x"f2",x"05",x"99"),
   670 => (x"01",x"ab",x"b7",x"c0"),
   671 => (x"c1",x"87",x"e1",x"fe"),
   672 => (x"f2",x"8e",x"f0",x"48"),
   673 => (x"5e",x"0e",x"87",x"c5"),
   674 => (x"0e",x"5d",x"5c",x"5b"),
   675 => (x"02",x"9b",x"4b",x"71"),
   676 => (x"a3",x"c8",x"87",x"c7"),
   677 => (x"c5",x"05",x"6d",x"4d"),
   678 => (x"c0",x"48",x"ff",x"87"),
   679 => (x"a3",x"d0",x"87",x"fd"),
   680 => (x"c7",x"49",x"6c",x"4c"),
   681 => (x"d8",x"05",x"99",x"ff"),
   682 => (x"c9",x"02",x"6c",x"87"),
   683 => (x"73",x"1e",x"c1",x"87"),
   684 => (x"87",x"ea",x"f6",x"49"),
   685 => (x"e5",x"c2",x"86",x"c4"),
   686 => (x"49",x"73",x"1e",x"e2"),
   687 => (x"c4",x"87",x"f9",x"f7"),
   688 => (x"6d",x"4a",x"6c",x"86"),
   689 => (x"87",x"c4",x"04",x"aa"),
   690 => (x"87",x"cf",x"48",x"ff"),
   691 => (x"72",x"7c",x"a2",x"c1"),
   692 => (x"99",x"ff",x"c7",x"49"),
   693 => (x"81",x"e2",x"e5",x"c2"),
   694 => (x"f0",x"48",x"69",x"97"),
   695 => (x"73",x"1e",x"87",x"ed"),
   696 => (x"9b",x"4b",x"71",x"1e"),
   697 => (x"87",x"e4",x"c0",x"02"),
   698 => (x"5b",x"cf",x"f2",x"c2"),
   699 => (x"8a",x"c2",x"4a",x"73"),
   700 => (x"bf",x"e2",x"ed",x"c2"),
   701 => (x"f1",x"c2",x"92",x"49"),
   702 => (x"72",x"48",x"bf",x"fb"),
   703 => (x"d3",x"f2",x"c2",x"80"),
   704 => (x"c4",x"48",x"71",x"58"),
   705 => (x"f2",x"ed",x"c2",x"30"),
   706 => (x"87",x"ed",x"c0",x"58"),
   707 => (x"48",x"cb",x"f2",x"c2"),
   708 => (x"bf",x"ff",x"f1",x"c2"),
   709 => (x"cf",x"f2",x"c2",x"78"),
   710 => (x"c3",x"f2",x"c2",x"48"),
   711 => (x"ed",x"c2",x"78",x"bf"),
   712 => (x"c9",x"02",x"bf",x"ea"),
   713 => (x"e2",x"ed",x"c2",x"87"),
   714 => (x"31",x"c4",x"49",x"bf"),
   715 => (x"f2",x"c2",x"87",x"c7"),
   716 => (x"c4",x"49",x"bf",x"c7"),
   717 => (x"f2",x"ed",x"c2",x"31"),
   718 => (x"87",x"d3",x"ef",x"59"),
   719 => (x"5c",x"5b",x"5e",x"0e"),
   720 => (x"c0",x"4a",x"71",x"0e"),
   721 => (x"02",x"9a",x"72",x"4b"),
   722 => (x"da",x"87",x"e1",x"c0"),
   723 => (x"69",x"9f",x"49",x"a2"),
   724 => (x"ea",x"ed",x"c2",x"4b"),
   725 => (x"87",x"cf",x"02",x"bf"),
   726 => (x"9f",x"49",x"a2",x"d4"),
   727 => (x"c0",x"4c",x"49",x"69"),
   728 => (x"d0",x"9c",x"ff",x"ff"),
   729 => (x"c0",x"87",x"c2",x"34"),
   730 => (x"b3",x"49",x"74",x"4c"),
   731 => (x"ed",x"fd",x"49",x"73"),
   732 => (x"87",x"d9",x"ee",x"87"),
   733 => (x"5c",x"5b",x"5e",x"0e"),
   734 => (x"86",x"f4",x"0e",x"5d"),
   735 => (x"7e",x"c0",x"4a",x"71"),
   736 => (x"d8",x"02",x"9a",x"72"),
   737 => (x"de",x"e5",x"c2",x"87"),
   738 => (x"c2",x"78",x"c0",x"48"),
   739 => (x"c2",x"48",x"d6",x"e5"),
   740 => (x"78",x"bf",x"cf",x"f2"),
   741 => (x"48",x"da",x"e5",x"c2"),
   742 => (x"bf",x"cb",x"f2",x"c2"),
   743 => (x"ff",x"ed",x"c2",x"78"),
   744 => (x"c2",x"50",x"c0",x"48"),
   745 => (x"49",x"bf",x"ee",x"ed"),
   746 => (x"bf",x"de",x"e5",x"c2"),
   747 => (x"03",x"aa",x"71",x"4a"),
   748 => (x"72",x"87",x"ca",x"c4"),
   749 => (x"05",x"99",x"cf",x"49"),
   750 => (x"c0",x"87",x"ea",x"c0"),
   751 => (x"c2",x"48",x"d0",x"f5"),
   752 => (x"78",x"bf",x"d6",x"e5"),
   753 => (x"1e",x"e2",x"e5",x"c2"),
   754 => (x"bf",x"d6",x"e5",x"c2"),
   755 => (x"d6",x"e5",x"c2",x"49"),
   756 => (x"78",x"a1",x"c1",x"48"),
   757 => (x"f4",x"de",x"ff",x"71"),
   758 => (x"c0",x"86",x"c4",x"87"),
   759 => (x"c2",x"48",x"cc",x"f5"),
   760 => (x"cc",x"78",x"e2",x"e5"),
   761 => (x"cc",x"f5",x"c0",x"87"),
   762 => (x"e0",x"c0",x"48",x"bf"),
   763 => (x"d0",x"f5",x"c0",x"80"),
   764 => (x"de",x"e5",x"c2",x"58"),
   765 => (x"80",x"c1",x"48",x"bf"),
   766 => (x"58",x"e2",x"e5",x"c2"),
   767 => (x"00",x"0d",x"4c",x"27"),
   768 => (x"bf",x"97",x"bf",x"00"),
   769 => (x"c2",x"02",x"9d",x"4d"),
   770 => (x"e5",x"c3",x"87",x"e3"),
   771 => (x"dc",x"c2",x"02",x"ad"),
   772 => (x"cc",x"f5",x"c0",x"87"),
   773 => (x"a3",x"cb",x"4b",x"bf"),
   774 => (x"cf",x"4c",x"11",x"49"),
   775 => (x"d2",x"c1",x"05",x"ac"),
   776 => (x"df",x"49",x"75",x"87"),
   777 => (x"cd",x"89",x"c1",x"99"),
   778 => (x"f2",x"ed",x"c2",x"91"),
   779 => (x"4a",x"a3",x"c1",x"81"),
   780 => (x"a3",x"c3",x"51",x"12"),
   781 => (x"c5",x"51",x"12",x"4a"),
   782 => (x"51",x"12",x"4a",x"a3"),
   783 => (x"12",x"4a",x"a3",x"c7"),
   784 => (x"4a",x"a3",x"c9",x"51"),
   785 => (x"a3",x"ce",x"51",x"12"),
   786 => (x"d0",x"51",x"12",x"4a"),
   787 => (x"51",x"12",x"4a",x"a3"),
   788 => (x"12",x"4a",x"a3",x"d2"),
   789 => (x"4a",x"a3",x"d4",x"51"),
   790 => (x"a3",x"d6",x"51",x"12"),
   791 => (x"d8",x"51",x"12",x"4a"),
   792 => (x"51",x"12",x"4a",x"a3"),
   793 => (x"12",x"4a",x"a3",x"dc"),
   794 => (x"4a",x"a3",x"de",x"51"),
   795 => (x"7e",x"c1",x"51",x"12"),
   796 => (x"74",x"87",x"fa",x"c0"),
   797 => (x"05",x"99",x"c8",x"49"),
   798 => (x"74",x"87",x"eb",x"c0"),
   799 => (x"05",x"99",x"d0",x"49"),
   800 => (x"66",x"dc",x"87",x"d1"),
   801 => (x"87",x"cb",x"c0",x"02"),
   802 => (x"66",x"dc",x"49",x"73"),
   803 => (x"02",x"98",x"70",x"0f"),
   804 => (x"6e",x"87",x"d3",x"c0"),
   805 => (x"87",x"c6",x"c0",x"05"),
   806 => (x"48",x"f2",x"ed",x"c2"),
   807 => (x"f5",x"c0",x"50",x"c0"),
   808 => (x"c2",x"48",x"bf",x"cc"),
   809 => (x"ed",x"c2",x"87",x"e1"),
   810 => (x"50",x"c0",x"48",x"ff"),
   811 => (x"ee",x"ed",x"c2",x"7e"),
   812 => (x"e5",x"c2",x"49",x"bf"),
   813 => (x"71",x"4a",x"bf",x"de"),
   814 => (x"f6",x"fb",x"04",x"aa"),
   815 => (x"cf",x"f2",x"c2",x"87"),
   816 => (x"c8",x"c0",x"05",x"bf"),
   817 => (x"ea",x"ed",x"c2",x"87"),
   818 => (x"f8",x"c1",x"02",x"bf"),
   819 => (x"da",x"e5",x"c2",x"87"),
   820 => (x"fe",x"e8",x"49",x"bf"),
   821 => (x"c2",x"49",x"70",x"87"),
   822 => (x"c4",x"59",x"de",x"e5"),
   823 => (x"e5",x"c2",x"48",x"a6"),
   824 => (x"c2",x"78",x"bf",x"da"),
   825 => (x"02",x"bf",x"ea",x"ed"),
   826 => (x"c4",x"87",x"d8",x"c0"),
   827 => (x"ff",x"cf",x"49",x"66"),
   828 => (x"99",x"f8",x"ff",x"ff"),
   829 => (x"c5",x"c0",x"02",x"a9"),
   830 => (x"c0",x"4c",x"c0",x"87"),
   831 => (x"4c",x"c1",x"87",x"e1"),
   832 => (x"c4",x"87",x"dc",x"c0"),
   833 => (x"ff",x"cf",x"49",x"66"),
   834 => (x"02",x"a9",x"99",x"f8"),
   835 => (x"c8",x"87",x"c8",x"c0"),
   836 => (x"78",x"c0",x"48",x"a6"),
   837 => (x"c8",x"87",x"c5",x"c0"),
   838 => (x"78",x"c1",x"48",x"a6"),
   839 => (x"74",x"4c",x"66",x"c8"),
   840 => (x"e0",x"c0",x"05",x"9c"),
   841 => (x"49",x"66",x"c4",x"87"),
   842 => (x"ed",x"c2",x"89",x"c2"),
   843 => (x"91",x"4a",x"bf",x"e2"),
   844 => (x"bf",x"fb",x"f1",x"c2"),
   845 => (x"d6",x"e5",x"c2",x"4a"),
   846 => (x"78",x"a1",x"72",x"48"),
   847 => (x"48",x"de",x"e5",x"c2"),
   848 => (x"de",x"f9",x"78",x"c0"),
   849 => (x"f4",x"48",x"c0",x"87"),
   850 => (x"87",x"ff",x"e6",x"8e"),
   851 => (x"00",x"00",x"00",x"00"),
   852 => (x"ff",x"ff",x"ff",x"ff"),
   853 => (x"00",x"00",x"0d",x"5c"),
   854 => (x"00",x"00",x"0d",x"65"),
   855 => (x"33",x"54",x"41",x"46"),
   856 => (x"20",x"20",x"20",x"32"),
   857 => (x"54",x"41",x"46",x"00"),
   858 => (x"20",x"20",x"36",x"31"),
   859 => (x"c2",x"1e",x"00",x"20"),
   860 => (x"48",x"bf",x"d4",x"f2"),
   861 => (x"c9",x"05",x"a8",x"dd"),
   862 => (x"dd",x"c2",x"c1",x"87"),
   863 => (x"4a",x"49",x"70",x"87"),
   864 => (x"d4",x"ff",x"87",x"c8"),
   865 => (x"78",x"ff",x"c3",x"48"),
   866 => (x"48",x"72",x"4a",x"68"),
   867 => (x"c2",x"1e",x"4f",x"26"),
   868 => (x"48",x"bf",x"d4",x"f2"),
   869 => (x"c6",x"05",x"a8",x"dd"),
   870 => (x"e9",x"c1",x"c1",x"87"),
   871 => (x"ff",x"87",x"d9",x"87"),
   872 => (x"ff",x"c3",x"48",x"d4"),
   873 => (x"48",x"d0",x"ff",x"78"),
   874 => (x"ff",x"78",x"e1",x"c0"),
   875 => (x"78",x"d4",x"48",x"d4"),
   876 => (x"48",x"d3",x"f2",x"c2"),
   877 => (x"50",x"bf",x"d4",x"ff"),
   878 => (x"ff",x"1e",x"4f",x"26"),
   879 => (x"e0",x"c0",x"48",x"d0"),
   880 => (x"1e",x"4f",x"26",x"78"),
   881 => (x"70",x"87",x"e7",x"fe"),
   882 => (x"c6",x"02",x"99",x"49"),
   883 => (x"a9",x"fb",x"c0",x"87"),
   884 => (x"71",x"87",x"f1",x"05"),
   885 => (x"0e",x"4f",x"26",x"48"),
   886 => (x"0e",x"5c",x"5b",x"5e"),
   887 => (x"4c",x"c0",x"4b",x"71"),
   888 => (x"70",x"87",x"cb",x"fe"),
   889 => (x"c0",x"02",x"99",x"49"),
   890 => (x"ec",x"c0",x"87",x"f9"),
   891 => (x"f2",x"c0",x"02",x"a9"),
   892 => (x"a9",x"fb",x"c0",x"87"),
   893 => (x"87",x"eb",x"c0",x"02"),
   894 => (x"ac",x"b7",x"66",x"cc"),
   895 => (x"d0",x"87",x"c7",x"03"),
   896 => (x"87",x"c2",x"02",x"66"),
   897 => (x"99",x"71",x"53",x"71"),
   898 => (x"c1",x"87",x"c2",x"02"),
   899 => (x"87",x"de",x"fd",x"84"),
   900 => (x"02",x"99",x"49",x"70"),
   901 => (x"ec",x"c0",x"87",x"cd"),
   902 => (x"87",x"c7",x"02",x"a9"),
   903 => (x"05",x"a9",x"fb",x"c0"),
   904 => (x"d0",x"87",x"d5",x"ff"),
   905 => (x"87",x"c3",x"02",x"66"),
   906 => (x"c0",x"7b",x"97",x"c0"),
   907 => (x"c4",x"05",x"a9",x"ec"),
   908 => (x"c5",x"4a",x"74",x"87"),
   909 => (x"c0",x"4a",x"74",x"87"),
   910 => (x"48",x"72",x"8a",x"0a"),
   911 => (x"4d",x"26",x"87",x"c2"),
   912 => (x"4b",x"26",x"4c",x"26"),
   913 => (x"fc",x"1e",x"4f",x"26"),
   914 => (x"49",x"70",x"87",x"e4"),
   915 => (x"a9",x"b7",x"f0",x"c0"),
   916 => (x"c0",x"87",x"ca",x"04"),
   917 => (x"01",x"a9",x"b7",x"f9"),
   918 => (x"f0",x"c0",x"87",x"c3"),
   919 => (x"b7",x"c1",x"c1",x"89"),
   920 => (x"87",x"ca",x"04",x"a9"),
   921 => (x"a9",x"b7",x"da",x"c1"),
   922 => (x"c0",x"87",x"c3",x"01"),
   923 => (x"48",x"71",x"89",x"f7"),
   924 => (x"5e",x"0e",x"4f",x"26"),
   925 => (x"71",x"0e",x"5c",x"5b"),
   926 => (x"4c",x"d4",x"ff",x"4a"),
   927 => (x"e9",x"c0",x"49",x"72"),
   928 => (x"9b",x"4b",x"70",x"87"),
   929 => (x"c1",x"87",x"c2",x"02"),
   930 => (x"48",x"d0",x"ff",x"8b"),
   931 => (x"d5",x"c1",x"78",x"c5"),
   932 => (x"c6",x"49",x"73",x"7c"),
   933 => (x"cc",x"e7",x"c1",x"31"),
   934 => (x"48",x"4a",x"bf",x"97"),
   935 => (x"7c",x"70",x"b0",x"71"),
   936 => (x"c4",x"48",x"d0",x"ff"),
   937 => (x"fe",x"48",x"73",x"78"),
   938 => (x"5e",x"0e",x"87",x"d6"),
   939 => (x"0e",x"5d",x"5c",x"5b"),
   940 => (x"4c",x"71",x"86",x"f4"),
   941 => (x"c0",x"48",x"a6",x"c4"),
   942 => (x"7e",x"a4",x"c8",x"78"),
   943 => (x"49",x"bf",x"97",x"6e"),
   944 => (x"05",x"a9",x"c1",x"c1"),
   945 => (x"a4",x"c9",x"87",x"dd"),
   946 => (x"49",x"69",x"97",x"49"),
   947 => (x"05",x"a9",x"d2",x"c1"),
   948 => (x"a4",x"ca",x"87",x"d1"),
   949 => (x"49",x"69",x"97",x"49"),
   950 => (x"05",x"a9",x"c3",x"c1"),
   951 => (x"48",x"df",x"87",x"c5"),
   952 => (x"fa",x"87",x"e1",x"c2"),
   953 => (x"4b",x"c0",x"87",x"e8"),
   954 => (x"97",x"c9",x"fe",x"c0"),
   955 => (x"a9",x"c0",x"49",x"bf"),
   956 => (x"fb",x"87",x"cf",x"04"),
   957 => (x"83",x"c1",x"87",x"cd"),
   958 => (x"97",x"c9",x"fe",x"c0"),
   959 => (x"06",x"ab",x"49",x"bf"),
   960 => (x"fe",x"c0",x"87",x"f1"),
   961 => (x"02",x"bf",x"97",x"c9"),
   962 => (x"e1",x"f9",x"87",x"cf"),
   963 => (x"99",x"49",x"70",x"87"),
   964 => (x"c0",x"87",x"c6",x"02"),
   965 => (x"f1",x"05",x"a9",x"ec"),
   966 => (x"f9",x"4b",x"c0",x"87"),
   967 => (x"4d",x"70",x"87",x"d0"),
   968 => (x"cc",x"87",x"cb",x"f9"),
   969 => (x"c5",x"f9",x"58",x"a6"),
   970 => (x"c1",x"4a",x"70",x"87"),
   971 => (x"bf",x"97",x"6e",x"83"),
   972 => (x"c7",x"02",x"ad",x"49"),
   973 => (x"ad",x"ff",x"c0",x"87"),
   974 => (x"87",x"ea",x"c0",x"05"),
   975 => (x"97",x"49",x"a4",x"c9"),
   976 => (x"66",x"c8",x"49",x"69"),
   977 => (x"87",x"c7",x"02",x"a9"),
   978 => (x"a8",x"ff",x"c0",x"48"),
   979 => (x"ca",x"87",x"d7",x"05"),
   980 => (x"69",x"97",x"49",x"a4"),
   981 => (x"c6",x"02",x"aa",x"49"),
   982 => (x"aa",x"ff",x"c0",x"87"),
   983 => (x"c4",x"87",x"c7",x"05"),
   984 => (x"78",x"c1",x"48",x"a6"),
   985 => (x"ec",x"c0",x"87",x"d3"),
   986 => (x"87",x"c6",x"02",x"ad"),
   987 => (x"05",x"ad",x"fb",x"c0"),
   988 => (x"4b",x"c0",x"87",x"c7"),
   989 => (x"c1",x"48",x"a6",x"c4"),
   990 => (x"02",x"66",x"c4",x"78"),
   991 => (x"f8",x"87",x"dc",x"fe"),
   992 => (x"48",x"73",x"87",x"f8"),
   993 => (x"f5",x"fa",x"8e",x"f4"),
   994 => (x"5e",x"0e",x"00",x"87"),
   995 => (x"0e",x"5d",x"5c",x"5b"),
   996 => (x"4d",x"71",x"86",x"f8"),
   997 => (x"75",x"4b",x"d4",x"ff"),
   998 => (x"d8",x"f2",x"c2",x"1e"),
   999 => (x"e4",x"df",x"ff",x"49"),
  1000 => (x"70",x"86",x"c4",x"87"),
  1001 => (x"fb",x"c4",x"02",x"98"),
  1002 => (x"ce",x"e7",x"c1",x"87"),
  1003 => (x"49",x"75",x"7e",x"bf"),
  1004 => (x"de",x"87",x"ff",x"fa"),
  1005 => (x"eb",x"c0",x"05",x"a8"),
  1006 => (x"c0",x"49",x"75",x"87"),
  1007 => (x"70",x"87",x"f9",x"f6"),
  1008 => (x"87",x"db",x"02",x"98"),
  1009 => (x"bf",x"fc",x"f6",x"c2"),
  1010 => (x"49",x"e1",x"c0",x"1e"),
  1011 => (x"87",x"c8",x"f4",x"c0"),
  1012 => (x"e7",x"c1",x"86",x"c4"),
  1013 => (x"50",x"c0",x"48",x"cc"),
  1014 => (x"49",x"c8",x"f7",x"c2"),
  1015 => (x"c1",x"87",x"eb",x"fe"),
  1016 => (x"87",x"c2",x"c4",x"48"),
  1017 => (x"c5",x"48",x"d0",x"ff"),
  1018 => (x"7b",x"d6",x"c1",x"78"),
  1019 => (x"a2",x"75",x"4a",x"c0"),
  1020 => (x"c1",x"7b",x"11",x"49"),
  1021 => (x"aa",x"b7",x"cb",x"82"),
  1022 => (x"cc",x"87",x"f3",x"04"),
  1023 => (x"7b",x"ff",x"c3",x"4a"),
  1024 => (x"e0",x"c0",x"82",x"c1"),
  1025 => (x"f4",x"04",x"aa",x"b7"),
  1026 => (x"48",x"d0",x"ff",x"87"),
  1027 => (x"ff",x"c3",x"78",x"c4"),
  1028 => (x"c1",x"78",x"c5",x"7b"),
  1029 => (x"7b",x"c1",x"7b",x"d3"),
  1030 => (x"48",x"6e",x"78",x"c4"),
  1031 => (x"06",x"a8",x"b7",x"c0"),
  1032 => (x"c2",x"87",x"f0",x"c2"),
  1033 => (x"4c",x"bf",x"e0",x"f2"),
  1034 => (x"88",x"74",x"48",x"6e"),
  1035 => (x"9c",x"74",x"7e",x"70"),
  1036 => (x"87",x"fd",x"c1",x"02"),
  1037 => (x"4d",x"e2",x"e5",x"c2"),
  1038 => (x"c8",x"48",x"a6",x"c4"),
  1039 => (x"c0",x"8c",x"78",x"c0"),
  1040 => (x"c6",x"03",x"ac",x"b7"),
  1041 => (x"a4",x"c0",x"c8",x"87"),
  1042 => (x"c2",x"4c",x"c0",x"78"),
  1043 => (x"bf",x"97",x"d3",x"f2"),
  1044 => (x"02",x"99",x"d0",x"49"),
  1045 => (x"1e",x"c0",x"87",x"d1"),
  1046 => (x"49",x"d8",x"f2",x"c2"),
  1047 => (x"c4",x"87",x"d9",x"e1"),
  1048 => (x"4a",x"49",x"70",x"86"),
  1049 => (x"c2",x"87",x"ee",x"c0"),
  1050 => (x"c2",x"1e",x"e2",x"e5"),
  1051 => (x"e1",x"49",x"d8",x"f2"),
  1052 => (x"86",x"c4",x"87",x"c6"),
  1053 => (x"ff",x"4a",x"49",x"70"),
  1054 => (x"c5",x"c8",x"48",x"d0"),
  1055 => (x"7b",x"d4",x"c1",x"78"),
  1056 => (x"66",x"c4",x"7b",x"15"),
  1057 => (x"c8",x"88",x"c1",x"48"),
  1058 => (x"98",x"70",x"58",x"a6"),
  1059 => (x"87",x"f0",x"ff",x"05"),
  1060 => (x"c4",x"48",x"d0",x"ff"),
  1061 => (x"05",x"9a",x"72",x"78"),
  1062 => (x"48",x"c0",x"87",x"c5"),
  1063 => (x"c1",x"87",x"c7",x"c1"),
  1064 => (x"d8",x"f2",x"c2",x"1e"),
  1065 => (x"f5",x"de",x"ff",x"49"),
  1066 => (x"74",x"86",x"c4",x"87"),
  1067 => (x"c3",x"fe",x"05",x"9c"),
  1068 => (x"c0",x"48",x"6e",x"87"),
  1069 => (x"d1",x"06",x"a8",x"b7"),
  1070 => (x"d8",x"f2",x"c2",x"87"),
  1071 => (x"d0",x"78",x"c0",x"48"),
  1072 => (x"f4",x"78",x"c0",x"80"),
  1073 => (x"e4",x"f2",x"c2",x"80"),
  1074 => (x"48",x"6e",x"78",x"bf"),
  1075 => (x"01",x"a8",x"b7",x"c0"),
  1076 => (x"ff",x"87",x"d0",x"fd"),
  1077 => (x"78",x"c5",x"48",x"d0"),
  1078 => (x"c0",x"7b",x"d3",x"c1"),
  1079 => (x"c1",x"78",x"c4",x"7b"),
  1080 => (x"87",x"c2",x"c0",x"48"),
  1081 => (x"8e",x"f8",x"48",x"c0"),
  1082 => (x"4c",x"26",x"4d",x"26"),
  1083 => (x"4f",x"26",x"4b",x"26"),
  1084 => (x"5c",x"5b",x"5e",x"0e"),
  1085 => (x"71",x"1e",x"0e",x"5d"),
  1086 => (x"4d",x"4c",x"c0",x"4b"),
  1087 => (x"e8",x"c0",x"04",x"ab"),
  1088 => (x"ea",x"fa",x"c0",x"87"),
  1089 => (x"02",x"9d",x"75",x"1e"),
  1090 => (x"4a",x"c0",x"87",x"c4"),
  1091 => (x"4a",x"c1",x"87",x"c2"),
  1092 => (x"df",x"e9",x"49",x"72"),
  1093 => (x"70",x"86",x"c4",x"87"),
  1094 => (x"6e",x"84",x"c1",x"7e"),
  1095 => (x"73",x"87",x"c2",x"05"),
  1096 => (x"73",x"85",x"c1",x"4c"),
  1097 => (x"d8",x"ff",x"06",x"ac"),
  1098 => (x"26",x"48",x"6e",x"87"),
  1099 => (x"1e",x"87",x"f9",x"fe"),
  1100 => (x"66",x"c4",x"4a",x"71"),
  1101 => (x"72",x"87",x"c5",x"05"),
  1102 => (x"87",x"ce",x"f9",x"49"),
  1103 => (x"5e",x"0e",x"4f",x"26"),
  1104 => (x"0e",x"5d",x"5c",x"5b"),
  1105 => (x"49",x"4c",x"71",x"1e"),
  1106 => (x"f3",x"c2",x"91",x"de"),
  1107 => (x"85",x"71",x"4d",x"c0"),
  1108 => (x"c1",x"02",x"6d",x"97"),
  1109 => (x"f2",x"c2",x"87",x"dc"),
  1110 => (x"74",x"4a",x"bf",x"ec"),
  1111 => (x"fe",x"49",x"72",x"82"),
  1112 => (x"7e",x"70",x"87",x"ce"),
  1113 => (x"f2",x"c0",x"02",x"6e"),
  1114 => (x"f4",x"f2",x"c2",x"87"),
  1115 => (x"cb",x"4a",x"6e",x"4b"),
  1116 => (x"f3",x"fc",x"fe",x"49"),
  1117 => (x"cb",x"4b",x"74",x"87"),
  1118 => (x"e0",x"e7",x"c1",x"93"),
  1119 => (x"c1",x"83",x"c4",x"83"),
  1120 => (x"74",x"7b",x"f6",x"c6"),
  1121 => (x"d0",x"cb",x"c1",x"49"),
  1122 => (x"c1",x"7b",x"75",x"87"),
  1123 => (x"bf",x"97",x"cd",x"e7"),
  1124 => (x"f2",x"c2",x"1e",x"49"),
  1125 => (x"d6",x"fe",x"49",x"f4"),
  1126 => (x"74",x"86",x"c4",x"87"),
  1127 => (x"f8",x"ca",x"c1",x"49"),
  1128 => (x"c1",x"49",x"c0",x"87"),
  1129 => (x"c2",x"87",x"d7",x"cc"),
  1130 => (x"c0",x"48",x"d4",x"f2"),
  1131 => (x"dd",x"49",x"c1",x"78"),
  1132 => (x"fc",x"26",x"87",x"d9"),
  1133 => (x"6f",x"4c",x"87",x"f2"),
  1134 => (x"6e",x"69",x"64",x"61"),
  1135 => (x"2e",x"2e",x"2e",x"67"),
  1136 => (x"5b",x"5e",x"0e",x"00"),
  1137 => (x"4b",x"71",x"0e",x"5c"),
  1138 => (x"ec",x"f2",x"c2",x"4a"),
  1139 => (x"49",x"72",x"82",x"bf"),
  1140 => (x"70",x"87",x"dd",x"fc"),
  1141 => (x"c4",x"02",x"9c",x"4c"),
  1142 => (x"df",x"e5",x"49",x"87"),
  1143 => (x"ec",x"f2",x"c2",x"87"),
  1144 => (x"c1",x"78",x"c0",x"48"),
  1145 => (x"87",x"e3",x"dc",x"49"),
  1146 => (x"0e",x"87",x"ff",x"fb"),
  1147 => (x"5d",x"5c",x"5b",x"5e"),
  1148 => (x"c2",x"86",x"f4",x"0e"),
  1149 => (x"c0",x"4d",x"e2",x"e5"),
  1150 => (x"48",x"a6",x"c4",x"4c"),
  1151 => (x"f2",x"c2",x"78",x"c0"),
  1152 => (x"c0",x"49",x"bf",x"ec"),
  1153 => (x"c1",x"c1",x"06",x"a9"),
  1154 => (x"e2",x"e5",x"c2",x"87"),
  1155 => (x"c0",x"02",x"98",x"48"),
  1156 => (x"fa",x"c0",x"87",x"f8"),
  1157 => (x"66",x"c8",x"1e",x"ea"),
  1158 => (x"c4",x"87",x"c7",x"02"),
  1159 => (x"78",x"c0",x"48",x"a6"),
  1160 => (x"a6",x"c4",x"87",x"c5"),
  1161 => (x"c4",x"78",x"c1",x"48"),
  1162 => (x"c7",x"e5",x"49",x"66"),
  1163 => (x"70",x"86",x"c4",x"87"),
  1164 => (x"c4",x"84",x"c1",x"4d"),
  1165 => (x"80",x"c1",x"48",x"66"),
  1166 => (x"c2",x"58",x"a6",x"c8"),
  1167 => (x"49",x"bf",x"ec",x"f2"),
  1168 => (x"87",x"c6",x"03",x"ac"),
  1169 => (x"ff",x"05",x"9d",x"75"),
  1170 => (x"4c",x"c0",x"87",x"c8"),
  1171 => (x"c3",x"02",x"9d",x"75"),
  1172 => (x"fa",x"c0",x"87",x"e0"),
  1173 => (x"66",x"c8",x"1e",x"ea"),
  1174 => (x"cc",x"87",x"c7",x"02"),
  1175 => (x"78",x"c0",x"48",x"a6"),
  1176 => (x"a6",x"cc",x"87",x"c5"),
  1177 => (x"cc",x"78",x"c1",x"48"),
  1178 => (x"c7",x"e4",x"49",x"66"),
  1179 => (x"70",x"86",x"c4",x"87"),
  1180 => (x"c2",x"02",x"6e",x"7e"),
  1181 => (x"49",x"6e",x"87",x"e9"),
  1182 => (x"69",x"97",x"81",x"cb"),
  1183 => (x"02",x"99",x"d0",x"49"),
  1184 => (x"c1",x"87",x"d6",x"c1"),
  1185 => (x"74",x"4a",x"c1",x"c7"),
  1186 => (x"c1",x"91",x"cb",x"49"),
  1187 => (x"72",x"81",x"e0",x"e7"),
  1188 => (x"c3",x"81",x"c8",x"79"),
  1189 => (x"49",x"74",x"51",x"ff"),
  1190 => (x"f3",x"c2",x"91",x"de"),
  1191 => (x"85",x"71",x"4d",x"c0"),
  1192 => (x"7d",x"97",x"c1",x"c2"),
  1193 => (x"c0",x"49",x"a5",x"c1"),
  1194 => (x"ed",x"c2",x"51",x"e0"),
  1195 => (x"02",x"bf",x"97",x"f2"),
  1196 => (x"84",x"c1",x"87",x"d2"),
  1197 => (x"c2",x"4b",x"a5",x"c2"),
  1198 => (x"db",x"4a",x"f2",x"ed"),
  1199 => (x"e7",x"f7",x"fe",x"49"),
  1200 => (x"87",x"db",x"c1",x"87"),
  1201 => (x"c0",x"49",x"a5",x"cd"),
  1202 => (x"c2",x"84",x"c1",x"51"),
  1203 => (x"4a",x"6e",x"4b",x"a5"),
  1204 => (x"f7",x"fe",x"49",x"cb"),
  1205 => (x"c6",x"c1",x"87",x"d2"),
  1206 => (x"fe",x"c4",x"c1",x"87"),
  1207 => (x"cb",x"49",x"74",x"4a"),
  1208 => (x"e0",x"e7",x"c1",x"91"),
  1209 => (x"c2",x"79",x"72",x"81"),
  1210 => (x"bf",x"97",x"f2",x"ed"),
  1211 => (x"74",x"87",x"d8",x"02"),
  1212 => (x"c1",x"91",x"de",x"49"),
  1213 => (x"c0",x"f3",x"c2",x"84"),
  1214 => (x"c2",x"83",x"71",x"4b"),
  1215 => (x"dd",x"4a",x"f2",x"ed"),
  1216 => (x"e3",x"f6",x"fe",x"49"),
  1217 => (x"74",x"87",x"d8",x"87"),
  1218 => (x"c2",x"93",x"de",x"4b"),
  1219 => (x"cb",x"83",x"c0",x"f3"),
  1220 => (x"51",x"c0",x"49",x"a3"),
  1221 => (x"6e",x"73",x"84",x"c1"),
  1222 => (x"fe",x"49",x"cb",x"4a"),
  1223 => (x"c4",x"87",x"c9",x"f6"),
  1224 => (x"80",x"c1",x"48",x"66"),
  1225 => (x"c7",x"58",x"a6",x"c8"),
  1226 => (x"c5",x"c0",x"03",x"ac"),
  1227 => (x"fc",x"05",x"6e",x"87"),
  1228 => (x"48",x"74",x"87",x"e0"),
  1229 => (x"ef",x"f6",x"8e",x"f4"),
  1230 => (x"1e",x"73",x"1e",x"87"),
  1231 => (x"cb",x"49",x"4b",x"71"),
  1232 => (x"e0",x"e7",x"c1",x"91"),
  1233 => (x"4a",x"a1",x"c8",x"81"),
  1234 => (x"48",x"cc",x"e7",x"c1"),
  1235 => (x"a1",x"c9",x"50",x"12"),
  1236 => (x"c9",x"fe",x"c0",x"4a"),
  1237 => (x"ca",x"50",x"12",x"48"),
  1238 => (x"cd",x"e7",x"c1",x"81"),
  1239 => (x"c1",x"50",x"11",x"48"),
  1240 => (x"bf",x"97",x"cd",x"e7"),
  1241 => (x"49",x"c0",x"1e",x"49"),
  1242 => (x"c2",x"87",x"c4",x"f7"),
  1243 => (x"de",x"48",x"d4",x"f2"),
  1244 => (x"d6",x"49",x"c1",x"78"),
  1245 => (x"f5",x"26",x"87",x"d5"),
  1246 => (x"71",x"1e",x"87",x"f2"),
  1247 => (x"91",x"cb",x"49",x"4a"),
  1248 => (x"81",x"e0",x"e7",x"c1"),
  1249 => (x"48",x"11",x"81",x"c8"),
  1250 => (x"58",x"d8",x"f2",x"c2"),
  1251 => (x"48",x"ec",x"f2",x"c2"),
  1252 => (x"49",x"c1",x"78",x"c0"),
  1253 => (x"26",x"87",x"f4",x"d5"),
  1254 => (x"49",x"c0",x"1e",x"4f"),
  1255 => (x"87",x"de",x"c4",x"c1"),
  1256 => (x"71",x"1e",x"4f",x"26"),
  1257 => (x"87",x"d2",x"02",x"99"),
  1258 => (x"48",x"f5",x"e8",x"c1"),
  1259 => (x"80",x"f7",x"50",x"c0"),
  1260 => (x"40",x"fa",x"cd",x"c1"),
  1261 => (x"78",x"d9",x"e7",x"c1"),
  1262 => (x"e8",x"c1",x"87",x"ce"),
  1263 => (x"e7",x"c1",x"48",x"f1"),
  1264 => (x"80",x"fc",x"78",x"d2"),
  1265 => (x"78",x"d9",x"ce",x"c1"),
  1266 => (x"5e",x"0e",x"4f",x"26"),
  1267 => (x"71",x"0e",x"5c",x"5b"),
  1268 => (x"92",x"cb",x"4a",x"4c"),
  1269 => (x"82",x"e0",x"e7",x"c1"),
  1270 => (x"c9",x"49",x"a2",x"c8"),
  1271 => (x"6b",x"97",x"4b",x"a2"),
  1272 => (x"69",x"97",x"1e",x"4b"),
  1273 => (x"82",x"ca",x"1e",x"49"),
  1274 => (x"e5",x"c0",x"49",x"12"),
  1275 => (x"49",x"c0",x"87",x"ca"),
  1276 => (x"74",x"87",x"d8",x"d4"),
  1277 => (x"e0",x"c1",x"c1",x"49"),
  1278 => (x"f3",x"8e",x"f8",x"87"),
  1279 => (x"73",x"1e",x"87",x"ec"),
  1280 => (x"49",x"4b",x"71",x"1e"),
  1281 => (x"73",x"87",x"c3",x"ff"),
  1282 => (x"87",x"fe",x"fe",x"49"),
  1283 => (x"1e",x"87",x"dd",x"f3"),
  1284 => (x"4b",x"71",x"1e",x"73"),
  1285 => (x"02",x"4a",x"a3",x"c6"),
  1286 => (x"8a",x"c1",x"87",x"db"),
  1287 => (x"8a",x"87",x"d6",x"02"),
  1288 => (x"87",x"da",x"c1",x"02"),
  1289 => (x"fc",x"c0",x"02",x"8a"),
  1290 => (x"c0",x"02",x"8a",x"87"),
  1291 => (x"02",x"8a",x"87",x"e1"),
  1292 => (x"db",x"c1",x"87",x"cb"),
  1293 => (x"fd",x"49",x"c7",x"87"),
  1294 => (x"de",x"c1",x"87",x"c0"),
  1295 => (x"ec",x"f2",x"c2",x"87"),
  1296 => (x"cb",x"c1",x"02",x"bf"),
  1297 => (x"88",x"c1",x"48",x"87"),
  1298 => (x"58",x"f0",x"f2",x"c2"),
  1299 => (x"c2",x"87",x"c1",x"c1"),
  1300 => (x"02",x"bf",x"f0",x"f2"),
  1301 => (x"c2",x"87",x"f9",x"c0"),
  1302 => (x"48",x"bf",x"ec",x"f2"),
  1303 => (x"f2",x"c2",x"80",x"c1"),
  1304 => (x"eb",x"c0",x"58",x"f0"),
  1305 => (x"ec",x"f2",x"c2",x"87"),
  1306 => (x"89",x"c6",x"49",x"bf"),
  1307 => (x"59",x"f0",x"f2",x"c2"),
  1308 => (x"03",x"a9",x"b7",x"c0"),
  1309 => (x"f2",x"c2",x"87",x"da"),
  1310 => (x"78",x"c0",x"48",x"ec"),
  1311 => (x"f2",x"c2",x"87",x"d2"),
  1312 => (x"cb",x"02",x"bf",x"f0"),
  1313 => (x"ec",x"f2",x"c2",x"87"),
  1314 => (x"80",x"c6",x"48",x"bf"),
  1315 => (x"58",x"f0",x"f2",x"c2"),
  1316 => (x"f6",x"d1",x"49",x"c0"),
  1317 => (x"c0",x"49",x"73",x"87"),
  1318 => (x"f1",x"87",x"fe",x"fe"),
  1319 => (x"73",x"1e",x"87",x"ce"),
  1320 => (x"c2",x"4b",x"71",x"1e"),
  1321 => (x"dd",x"48",x"d4",x"f2"),
  1322 => (x"d1",x"49",x"c0",x"78"),
  1323 => (x"49",x"73",x"87",x"dd"),
  1324 => (x"87",x"e5",x"fe",x"c0"),
  1325 => (x"0e",x"87",x"f5",x"f0"),
  1326 => (x"5d",x"5c",x"5b",x"5e"),
  1327 => (x"86",x"cc",x"ff",x"0e"),
  1328 => (x"c8",x"59",x"a6",x"d8"),
  1329 => (x"78",x"c0",x"48",x"a6"),
  1330 => (x"c8",x"c1",x"80",x"c4"),
  1331 => (x"80",x"c4",x"78",x"66"),
  1332 => (x"f2",x"c2",x"78",x"c1"),
  1333 => (x"78",x"c1",x"48",x"f0"),
  1334 => (x"bf",x"d4",x"f2",x"c2"),
  1335 => (x"05",x"a8",x"de",x"48"),
  1336 => (x"c6",x"f4",x"87",x"cb"),
  1337 => (x"cc",x"49",x"70",x"87"),
  1338 => (x"d0",x"cf",x"59",x"a6"),
  1339 => (x"87",x"de",x"e2",x"87"),
  1340 => (x"e1",x"87",x"d0",x"e3"),
  1341 => (x"4c",x"70",x"87",x"f8"),
  1342 => (x"c1",x"05",x"66",x"d4"),
  1343 => (x"c4",x"c1",x"87",x"fc"),
  1344 => (x"80",x"c4",x"48",x"66"),
  1345 => (x"a6",x"c4",x"7e",x"70"),
  1346 => (x"78",x"bf",x"6e",x"48"),
  1347 => (x"e3",x"c1",x"1e",x"72"),
  1348 => (x"66",x"c8",x"48",x"f2"),
  1349 => (x"4a",x"a1",x"c8",x"49"),
  1350 => (x"aa",x"71",x"41",x"20"),
  1351 => (x"10",x"87",x"f9",x"05"),
  1352 => (x"c1",x"4a",x"26",x"51"),
  1353 => (x"c1",x"48",x"66",x"c4"),
  1354 => (x"6e",x"78",x"f9",x"cc"),
  1355 => (x"81",x"c7",x"49",x"bf"),
  1356 => (x"c4",x"c1",x"51",x"74"),
  1357 => (x"81",x"c8",x"49",x"66"),
  1358 => (x"c4",x"c1",x"51",x"c1"),
  1359 => (x"81",x"c9",x"49",x"66"),
  1360 => (x"c4",x"c1",x"51",x"c0"),
  1361 => (x"81",x"ca",x"49",x"66"),
  1362 => (x"fb",x"c0",x"51",x"c0"),
  1363 => (x"87",x"cf",x"02",x"ac"),
  1364 => (x"1e",x"d8",x"1e",x"c1"),
  1365 => (x"49",x"bf",x"66",x"c8"),
  1366 => (x"fa",x"e1",x"81",x"c8"),
  1367 => (x"c1",x"86",x"c8",x"87"),
  1368 => (x"c0",x"48",x"66",x"c8"),
  1369 => (x"87",x"c7",x"01",x"a8"),
  1370 => (x"c1",x"48",x"a6",x"c8"),
  1371 => (x"c1",x"87",x"ce",x"78"),
  1372 => (x"c1",x"48",x"66",x"c8"),
  1373 => (x"58",x"a6",x"d0",x"88"),
  1374 => (x"c6",x"e1",x"87",x"c3"),
  1375 => (x"48",x"a6",x"d8",x"87"),
  1376 => (x"9c",x"74",x"78",x"c2"),
  1377 => (x"87",x"f1",x"cc",x"02"),
  1378 => (x"c1",x"48",x"66",x"c8"),
  1379 => (x"03",x"a8",x"66",x"cc"),
  1380 => (x"dc",x"87",x"e6",x"cc"),
  1381 => (x"78",x"c0",x"48",x"a6"),
  1382 => (x"78",x"c0",x"80",x"c4"),
  1383 => (x"87",x"ce",x"df",x"ff"),
  1384 => (x"66",x"d4",x"4c",x"70"),
  1385 => (x"05",x"a8",x"dd",x"48"),
  1386 => (x"e0",x"c0",x"87",x"c7"),
  1387 => (x"66",x"d4",x"48",x"a6"),
  1388 => (x"ac",x"d0",x"c1",x"78"),
  1389 => (x"87",x"eb",x"c0",x"05"),
  1390 => (x"87",x"f2",x"de",x"ff"),
  1391 => (x"87",x"ee",x"de",x"ff"),
  1392 => (x"ec",x"c0",x"4c",x"70"),
  1393 => (x"87",x"c6",x"05",x"ac"),
  1394 => (x"87",x"f7",x"df",x"ff"),
  1395 => (x"d0",x"c1",x"4c",x"70"),
  1396 => (x"87",x"c8",x"05",x"ac"),
  1397 => (x"c1",x"48",x"66",x"d0"),
  1398 => (x"58",x"a6",x"d4",x"80"),
  1399 => (x"02",x"ac",x"d0",x"c1"),
  1400 => (x"c0",x"87",x"d5",x"ff"),
  1401 => (x"d4",x"48",x"a6",x"e4"),
  1402 => (x"e0",x"c0",x"78",x"66"),
  1403 => (x"e4",x"c0",x"48",x"66"),
  1404 => (x"ca",x"05",x"a8",x"66"),
  1405 => (x"e8",x"c0",x"87",x"d5"),
  1406 => (x"78",x"c0",x"48",x"a6"),
  1407 => (x"c0",x"80",x"dc",x"ff"),
  1408 => (x"c0",x"4d",x"74",x"78"),
  1409 => (x"c9",x"02",x"8d",x"fb"),
  1410 => (x"8d",x"c9",x"87",x"db"),
  1411 => (x"c2",x"87",x"db",x"02"),
  1412 => (x"f7",x"c1",x"02",x"8d"),
  1413 => (x"02",x"8d",x"c9",x"87"),
  1414 => (x"c4",x"87",x"d8",x"c4"),
  1415 => (x"c1",x"c1",x"02",x"8d"),
  1416 => (x"02",x"8d",x"c1",x"87"),
  1417 => (x"c8",x"87",x"cc",x"c4"),
  1418 => (x"66",x"c8",x"87",x"f5"),
  1419 => (x"c1",x"91",x"cb",x"49"),
  1420 => (x"c4",x"81",x"66",x"c4"),
  1421 => (x"7e",x"6a",x"4a",x"a1"),
  1422 => (x"e3",x"c1",x"1e",x"71"),
  1423 => (x"66",x"c4",x"48",x"fe"),
  1424 => (x"4a",x"a1",x"cc",x"49"),
  1425 => (x"aa",x"71",x"41",x"20"),
  1426 => (x"87",x"f8",x"ff",x"05"),
  1427 => (x"49",x"26",x"51",x"10"),
  1428 => (x"79",x"de",x"d2",x"c1"),
  1429 => (x"87",x"d6",x"dc",x"ff"),
  1430 => (x"a6",x"c4",x"4c",x"70"),
  1431 => (x"c8",x"78",x"c1",x"48"),
  1432 => (x"a6",x"dc",x"87",x"c3"),
  1433 => (x"78",x"f0",x"c0",x"48"),
  1434 => (x"87",x"c2",x"dc",x"ff"),
  1435 => (x"ec",x"c0",x"4c",x"70"),
  1436 => (x"c4",x"c0",x"02",x"ac"),
  1437 => (x"a6",x"e0",x"c0",x"87"),
  1438 => (x"ac",x"ec",x"c0",x"5c"),
  1439 => (x"ff",x"87",x"cd",x"02"),
  1440 => (x"70",x"87",x"eb",x"db"),
  1441 => (x"ac",x"ec",x"c0",x"4c"),
  1442 => (x"87",x"f3",x"ff",x"05"),
  1443 => (x"02",x"ac",x"ec",x"c0"),
  1444 => (x"ff",x"87",x"c4",x"c0"),
  1445 => (x"c0",x"87",x"d7",x"db"),
  1446 => (x"d0",x"1e",x"ca",x"1e"),
  1447 => (x"91",x"cb",x"49",x"66"),
  1448 => (x"48",x"66",x"cc",x"c1"),
  1449 => (x"a6",x"cc",x"80",x"71"),
  1450 => (x"48",x"66",x"c8",x"58"),
  1451 => (x"a6",x"d0",x"80",x"c4"),
  1452 => (x"bf",x"66",x"cc",x"58"),
  1453 => (x"de",x"dc",x"ff",x"49"),
  1454 => (x"de",x"1e",x"c1",x"87"),
  1455 => (x"bf",x"66",x"d4",x"1e"),
  1456 => (x"d2",x"dc",x"ff",x"49"),
  1457 => (x"70",x"86",x"d0",x"87"),
  1458 => (x"89",x"09",x"c0",x"49"),
  1459 => (x"59",x"a6",x"f0",x"c0"),
  1460 => (x"48",x"66",x"ec",x"c0"),
  1461 => (x"c0",x"06",x"a8",x"c0"),
  1462 => (x"ec",x"c0",x"87",x"ee"),
  1463 => (x"a8",x"dd",x"48",x"66"),
  1464 => (x"87",x"e4",x"c0",x"03"),
  1465 => (x"49",x"bf",x"66",x"c4"),
  1466 => (x"81",x"66",x"ec",x"c0"),
  1467 => (x"c0",x"51",x"e0",x"c0"),
  1468 => (x"c1",x"49",x"66",x"ec"),
  1469 => (x"bf",x"66",x"c4",x"81"),
  1470 => (x"51",x"c1",x"c2",x"81"),
  1471 => (x"49",x"66",x"ec",x"c0"),
  1472 => (x"66",x"c4",x"81",x"c2"),
  1473 => (x"51",x"c0",x"81",x"bf"),
  1474 => (x"cc",x"c1",x"48",x"6e"),
  1475 => (x"49",x"6e",x"78",x"f9"),
  1476 => (x"66",x"d8",x"81",x"c8"),
  1477 => (x"c9",x"49",x"6e",x"51"),
  1478 => (x"51",x"66",x"d0",x"81"),
  1479 => (x"81",x"ca",x"49",x"6e"),
  1480 => (x"d8",x"51",x"66",x"dc"),
  1481 => (x"80",x"c1",x"48",x"66"),
  1482 => (x"48",x"58",x"a6",x"dc"),
  1483 => (x"78",x"c1",x"80",x"ec"),
  1484 => (x"ff",x"87",x"f2",x"c4"),
  1485 => (x"70",x"87",x"cf",x"dc"),
  1486 => (x"a6",x"f0",x"c0",x"49"),
  1487 => (x"c5",x"dc",x"ff",x"59"),
  1488 => (x"c0",x"49",x"70",x"87"),
  1489 => (x"dc",x"59",x"a6",x"e0"),
  1490 => (x"ec",x"c0",x"48",x"66"),
  1491 => (x"ca",x"c0",x"05",x"a8"),
  1492 => (x"48",x"a6",x"dc",x"87"),
  1493 => (x"78",x"66",x"ec",x"c0"),
  1494 => (x"ff",x"87",x"c4",x"c0"),
  1495 => (x"c8",x"87",x"cf",x"d8"),
  1496 => (x"91",x"cb",x"49",x"66"),
  1497 => (x"48",x"66",x"c4",x"c1"),
  1498 => (x"7e",x"70",x"80",x"71"),
  1499 => (x"82",x"c8",x"4a",x"6e"),
  1500 => (x"81",x"ca",x"49",x"6e"),
  1501 => (x"51",x"66",x"ec",x"c0"),
  1502 => (x"c1",x"49",x"66",x"dc"),
  1503 => (x"66",x"ec",x"c0",x"81"),
  1504 => (x"71",x"48",x"c1",x"89"),
  1505 => (x"c1",x"49",x"70",x"30"),
  1506 => (x"7a",x"97",x"71",x"89"),
  1507 => (x"bf",x"dc",x"f6",x"c2"),
  1508 => (x"66",x"ec",x"c0",x"49"),
  1509 => (x"4a",x"6a",x"97",x"29"),
  1510 => (x"c0",x"98",x"71",x"48"),
  1511 => (x"6e",x"58",x"a6",x"f4"),
  1512 => (x"a6",x"81",x"c4",x"49"),
  1513 => (x"c0",x"78",x"69",x"48"),
  1514 => (x"c0",x"48",x"66",x"e4"),
  1515 => (x"02",x"a8",x"66",x"e0"),
  1516 => (x"dc",x"87",x"c8",x"c0"),
  1517 => (x"78",x"c0",x"48",x"a6"),
  1518 => (x"dc",x"87",x"c5",x"c0"),
  1519 => (x"78",x"c1",x"48",x"a6"),
  1520 => (x"c0",x"1e",x"66",x"dc"),
  1521 => (x"66",x"cc",x"1e",x"e0"),
  1522 => (x"ca",x"d8",x"ff",x"49"),
  1523 => (x"70",x"86",x"c8",x"87"),
  1524 => (x"ac",x"b7",x"c0",x"4c"),
  1525 => (x"87",x"db",x"c1",x"06"),
  1526 => (x"74",x"48",x"66",x"c4"),
  1527 => (x"58",x"a6",x"c8",x"80"),
  1528 => (x"74",x"49",x"e0",x"c0"),
  1529 => (x"4b",x"66",x"c4",x"89"),
  1530 => (x"4a",x"fb",x"e3",x"c1"),
  1531 => (x"f7",x"e2",x"fe",x"71"),
  1532 => (x"48",x"66",x"c4",x"87"),
  1533 => (x"a6",x"c8",x"80",x"c2"),
  1534 => (x"66",x"e8",x"c0",x"58"),
  1535 => (x"c0",x"80",x"c1",x"48"),
  1536 => (x"c0",x"58",x"a6",x"ec"),
  1537 => (x"c1",x"49",x"66",x"f0"),
  1538 => (x"02",x"a9",x"70",x"81"),
  1539 => (x"c0",x"87",x"c5",x"c0"),
  1540 => (x"87",x"c2",x"c0",x"4d"),
  1541 => (x"1e",x"75",x"4d",x"c1"),
  1542 => (x"c0",x"49",x"a4",x"c2"),
  1543 => (x"88",x"71",x"48",x"e0"),
  1544 => (x"cc",x"1e",x"49",x"70"),
  1545 => (x"d6",x"ff",x"49",x"66"),
  1546 => (x"86",x"c8",x"87",x"ed"),
  1547 => (x"01",x"a8",x"b7",x"c0"),
  1548 => (x"c0",x"87",x"c6",x"ff"),
  1549 => (x"c0",x"02",x"66",x"e8"),
  1550 => (x"49",x"6e",x"87",x"d1"),
  1551 => (x"e8",x"c0",x"81",x"c9"),
  1552 => (x"48",x"6e",x"51",x"66"),
  1553 => (x"78",x"ca",x"cf",x"c1"),
  1554 => (x"6e",x"87",x"cc",x"c0"),
  1555 => (x"c2",x"81",x"c9",x"49"),
  1556 => (x"c1",x"48",x"6e",x"51"),
  1557 => (x"c4",x"78",x"fe",x"cf"),
  1558 => (x"78",x"c1",x"48",x"a6"),
  1559 => (x"ff",x"87",x"c6",x"c0"),
  1560 => (x"70",x"87",x"e0",x"d5"),
  1561 => (x"02",x"66",x"c4",x"4c"),
  1562 => (x"c8",x"87",x"f5",x"c0"),
  1563 => (x"66",x"cc",x"48",x"66"),
  1564 => (x"cb",x"c0",x"04",x"a8"),
  1565 => (x"48",x"66",x"c8",x"87"),
  1566 => (x"a6",x"cc",x"80",x"c1"),
  1567 => (x"87",x"e0",x"c0",x"58"),
  1568 => (x"c1",x"48",x"66",x"cc"),
  1569 => (x"58",x"a6",x"d0",x"88"),
  1570 => (x"c1",x"87",x"d5",x"c0"),
  1571 => (x"c0",x"05",x"ac",x"c6"),
  1572 => (x"66",x"d8",x"87",x"c8"),
  1573 => (x"dc",x"80",x"c1",x"48"),
  1574 => (x"d4",x"ff",x"58",x"a6"),
  1575 => (x"4c",x"70",x"87",x"e5"),
  1576 => (x"c1",x"48",x"66",x"d0"),
  1577 => (x"58",x"a6",x"d4",x"80"),
  1578 => (x"c0",x"02",x"9c",x"74"),
  1579 => (x"66",x"c8",x"87",x"cb"),
  1580 => (x"66",x"cc",x"c1",x"48"),
  1581 => (x"da",x"f3",x"04",x"a8"),
  1582 => (x"fd",x"d3",x"ff",x"87"),
  1583 => (x"48",x"66",x"c8",x"87"),
  1584 => (x"c0",x"03",x"a8",x"c7"),
  1585 => (x"f2",x"c2",x"87",x"e5"),
  1586 => (x"78",x"c0",x"48",x"f0"),
  1587 => (x"cb",x"49",x"66",x"c8"),
  1588 => (x"66",x"c4",x"c1",x"91"),
  1589 => (x"4a",x"a1",x"c4",x"81"),
  1590 => (x"52",x"c0",x"4a",x"6a"),
  1591 => (x"48",x"66",x"c8",x"79"),
  1592 => (x"a6",x"cc",x"80",x"c1"),
  1593 => (x"04",x"a8",x"c7",x"58"),
  1594 => (x"ff",x"87",x"db",x"ff"),
  1595 => (x"df",x"ff",x"8e",x"cc"),
  1596 => (x"6f",x"4c",x"87",x"f6"),
  1597 => (x"2a",x"20",x"64",x"61"),
  1598 => (x"3a",x"00",x"20",x"2e"),
  1599 => (x"49",x"44",x"00",x"20"),
  1600 => (x"77",x"53",x"20",x"50"),
  1601 => (x"68",x"63",x"74",x"69"),
  1602 => (x"1e",x"00",x"73",x"65"),
  1603 => (x"4b",x"71",x"1e",x"73"),
  1604 => (x"87",x"c6",x"02",x"9b"),
  1605 => (x"48",x"ec",x"f2",x"c2"),
  1606 => (x"1e",x"c7",x"78",x"c0"),
  1607 => (x"bf",x"ec",x"f2",x"c2"),
  1608 => (x"e7",x"c1",x"1e",x"49"),
  1609 => (x"f2",x"c2",x"1e",x"e0"),
  1610 => (x"ee",x"49",x"bf",x"d4"),
  1611 => (x"86",x"cc",x"87",x"c9"),
  1612 => (x"bf",x"d4",x"f2",x"c2"),
  1613 => (x"87",x"ea",x"e9",x"49"),
  1614 => (x"c8",x"02",x"9b",x"73"),
  1615 => (x"e0",x"e7",x"c1",x"87"),
  1616 => (x"e6",x"ed",x"c0",x"49"),
  1617 => (x"e3",x"de",x"ff",x"87"),
  1618 => (x"cd",x"c7",x"1e",x"87"),
  1619 => (x"fe",x"49",x"c1",x"87"),
  1620 => (x"e5",x"fe",x"87",x"f9"),
  1621 => (x"98",x"70",x"87",x"e0"),
  1622 => (x"fe",x"87",x"cd",x"02"),
  1623 => (x"70",x"87",x"f9",x"ec"),
  1624 => (x"87",x"c4",x"02",x"98"),
  1625 => (x"87",x"c2",x"4a",x"c1"),
  1626 => (x"9a",x"72",x"4a",x"c0"),
  1627 => (x"c0",x"87",x"ce",x"05"),
  1628 => (x"de",x"e6",x"c1",x"1e"),
  1629 => (x"d0",x"f9",x"c0",x"49"),
  1630 => (x"fe",x"86",x"c4",x"87"),
  1631 => (x"f3",x"fb",x"c0",x"87"),
  1632 => (x"c1",x"1e",x"c0",x"87"),
  1633 => (x"c0",x"49",x"e9",x"e6"),
  1634 => (x"c0",x"87",x"fe",x"f8"),
  1635 => (x"f9",x"fd",x"c0",x"1e"),
  1636 => (x"c0",x"49",x"70",x"87"),
  1637 => (x"c2",x"87",x"f2",x"f8"),
  1638 => (x"8e",x"f8",x"87",x"ff"),
  1639 => (x"44",x"53",x"4f",x"26"),
  1640 => (x"69",x"61",x"66",x"20"),
  1641 => (x"2e",x"64",x"65",x"6c"),
  1642 => (x"6f",x"6f",x"42",x"00"),
  1643 => (x"67",x"6e",x"69",x"74"),
  1644 => (x"00",x"2e",x"2e",x"2e"),
  1645 => (x"ec",x"f2",x"c2",x"1e"),
  1646 => (x"c2",x"78",x"c0",x"48"),
  1647 => (x"c0",x"48",x"d4",x"f2"),
  1648 => (x"87",x"c5",x"fe",x"78"),
  1649 => (x"87",x"e1",x"fd",x"c0"),
  1650 => (x"4f",x"26",x"48",x"c0"),
  1651 => (x"00",x"01",x"00",x"00"),
  1652 => (x"20",x"80",x"00",x"00"),
  1653 => (x"74",x"69",x"78",x"45"),
  1654 => (x"42",x"20",x"80",x"00"),
  1655 => (x"00",x"6b",x"63",x"61"),
  1656 => (x"00",x"00",x"13",x"7a"),
  1657 => (x"00",x"00",x"2c",x"c0"),
  1658 => (x"7a",x"00",x"00",x"00"),
  1659 => (x"de",x"00",x"00",x"13"),
  1660 => (x"00",x"00",x"00",x"2c"),
  1661 => (x"13",x"7a",x"00",x"00"),
  1662 => (x"2c",x"fc",x"00",x"00"),
  1663 => (x"00",x"00",x"00",x"00"),
  1664 => (x"00",x"13",x"7a",x"00"),
  1665 => (x"00",x"2d",x"1a",x"00"),
  1666 => (x"00",x"00",x"00",x"00"),
  1667 => (x"00",x"00",x"13",x"7a"),
  1668 => (x"00",x"00",x"2d",x"38"),
  1669 => (x"7a",x"00",x"00",x"00"),
  1670 => (x"56",x"00",x"00",x"13"),
  1671 => (x"00",x"00",x"00",x"2d"),
  1672 => (x"13",x"7a",x"00",x"00"),
  1673 => (x"2d",x"74",x"00",x"00"),
  1674 => (x"00",x"00",x"00",x"00"),
  1675 => (x"00",x"13",x"7a",x"00"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"00",x"00",x"00",x"00"),
  1678 => (x"00",x"00",x"14",x"0f"),
  1679 => (x"00",x"00",x"00",x"00"),
  1680 => (x"1e",x"00",x"00",x"00"),
  1681 => (x"c0",x"48",x"f0",x"fe"),
  1682 => (x"79",x"09",x"cd",x"78"),
  1683 => (x"1e",x"4f",x"26",x"09"),
  1684 => (x"bf",x"f0",x"fe",x"1e"),
  1685 => (x"26",x"26",x"48",x"7e"),
  1686 => (x"f0",x"fe",x"1e",x"4f"),
  1687 => (x"26",x"78",x"c1",x"48"),
  1688 => (x"f0",x"fe",x"1e",x"4f"),
  1689 => (x"26",x"78",x"c0",x"48"),
  1690 => (x"4a",x"71",x"1e",x"4f"),
  1691 => (x"26",x"52",x"52",x"c0"),
  1692 => (x"5b",x"5e",x"0e",x"4f"),
  1693 => (x"f4",x"0e",x"5d",x"5c"),
  1694 => (x"97",x"4d",x"71",x"86"),
  1695 => (x"a5",x"c1",x"7e",x"6d"),
  1696 => (x"48",x"6c",x"97",x"4c"),
  1697 => (x"6e",x"58",x"a6",x"c8"),
  1698 => (x"a8",x"66",x"c4",x"48"),
  1699 => (x"ff",x"87",x"c5",x"05"),
  1700 => (x"87",x"e6",x"c0",x"48"),
  1701 => (x"c2",x"87",x"ca",x"ff"),
  1702 => (x"6c",x"97",x"49",x"a5"),
  1703 => (x"4b",x"a3",x"71",x"4b"),
  1704 => (x"97",x"4b",x"6b",x"97"),
  1705 => (x"48",x"6e",x"7e",x"6c"),
  1706 => (x"a6",x"c8",x"80",x"c1"),
  1707 => (x"cc",x"98",x"c7",x"58"),
  1708 => (x"97",x"70",x"58",x"a6"),
  1709 => (x"87",x"e1",x"fe",x"7c"),
  1710 => (x"8e",x"f4",x"48",x"73"),
  1711 => (x"4c",x"26",x"4d",x"26"),
  1712 => (x"4f",x"26",x"4b",x"26"),
  1713 => (x"5c",x"5b",x"5e",x"0e"),
  1714 => (x"71",x"86",x"f4",x"0e"),
  1715 => (x"4a",x"66",x"d8",x"4c"),
  1716 => (x"c2",x"9a",x"ff",x"c3"),
  1717 => (x"6c",x"97",x"4b",x"a4"),
  1718 => (x"49",x"a1",x"73",x"49"),
  1719 => (x"6c",x"97",x"51",x"72"),
  1720 => (x"c1",x"48",x"6e",x"7e"),
  1721 => (x"58",x"a6",x"c8",x"80"),
  1722 => (x"a6",x"cc",x"98",x"c7"),
  1723 => (x"f4",x"54",x"70",x"58"),
  1724 => (x"87",x"ca",x"ff",x"8e"),
  1725 => (x"e8",x"fd",x"1e",x"1e"),
  1726 => (x"4a",x"bf",x"e0",x"87"),
  1727 => (x"c0",x"e0",x"c0",x"49"),
  1728 => (x"87",x"cb",x"02",x"99"),
  1729 => (x"f6",x"c2",x"1e",x"72"),
  1730 => (x"f7",x"fe",x"49",x"d2"),
  1731 => (x"fc",x"86",x"c4",x"87"),
  1732 => (x"7e",x"70",x"87",x"fd"),
  1733 => (x"26",x"87",x"c2",x"fd"),
  1734 => (x"c2",x"1e",x"4f",x"26"),
  1735 => (x"fd",x"49",x"d2",x"f6"),
  1736 => (x"eb",x"c1",x"87",x"c7"),
  1737 => (x"da",x"fc",x"49",x"f4"),
  1738 => (x"87",x"c7",x"c4",x"87"),
  1739 => (x"ff",x"1e",x"4f",x"26"),
  1740 => (x"e1",x"c8",x"48",x"d0"),
  1741 => (x"48",x"d4",x"ff",x"78"),
  1742 => (x"66",x"c4",x"78",x"c5"),
  1743 => (x"c3",x"87",x"c3",x"02"),
  1744 => (x"66",x"c8",x"78",x"e0"),
  1745 => (x"ff",x"87",x"c6",x"02"),
  1746 => (x"f0",x"c3",x"48",x"d4"),
  1747 => (x"48",x"d4",x"ff",x"78"),
  1748 => (x"d0",x"ff",x"78",x"71"),
  1749 => (x"78",x"e1",x"c8",x"48"),
  1750 => (x"26",x"78",x"e0",x"c0"),
  1751 => (x"5b",x"5e",x"0e",x"4f"),
  1752 => (x"4c",x"71",x"0e",x"5c"),
  1753 => (x"49",x"d2",x"f6",x"c2"),
  1754 => (x"70",x"87",x"c6",x"fc"),
  1755 => (x"aa",x"b7",x"c0",x"4a"),
  1756 => (x"87",x"e2",x"c2",x"04"),
  1757 => (x"05",x"aa",x"f0",x"c3"),
  1758 => (x"f0",x"c1",x"87",x"c9"),
  1759 => (x"78",x"c1",x"48",x"e2"),
  1760 => (x"c3",x"87",x"c3",x"c2"),
  1761 => (x"c9",x"05",x"aa",x"e0"),
  1762 => (x"e6",x"f0",x"c1",x"87"),
  1763 => (x"c1",x"78",x"c1",x"48"),
  1764 => (x"f0",x"c1",x"87",x"f4"),
  1765 => (x"c6",x"02",x"bf",x"e6"),
  1766 => (x"a2",x"c0",x"c2",x"87"),
  1767 => (x"72",x"87",x"c2",x"4b"),
  1768 => (x"05",x"9c",x"74",x"4b"),
  1769 => (x"f0",x"c1",x"87",x"d1"),
  1770 => (x"c1",x"1e",x"bf",x"e2"),
  1771 => (x"1e",x"bf",x"e6",x"f0"),
  1772 => (x"f9",x"fd",x"49",x"72"),
  1773 => (x"c1",x"86",x"c8",x"87"),
  1774 => (x"02",x"bf",x"e2",x"f0"),
  1775 => (x"73",x"87",x"e0",x"c0"),
  1776 => (x"29",x"b7",x"c4",x"49"),
  1777 => (x"c2",x"f2",x"c1",x"91"),
  1778 => (x"cf",x"4a",x"73",x"81"),
  1779 => (x"c1",x"92",x"c2",x"9a"),
  1780 => (x"70",x"30",x"72",x"48"),
  1781 => (x"72",x"ba",x"ff",x"4a"),
  1782 => (x"70",x"98",x"69",x"48"),
  1783 => (x"73",x"87",x"db",x"79"),
  1784 => (x"29",x"b7",x"c4",x"49"),
  1785 => (x"c2",x"f2",x"c1",x"91"),
  1786 => (x"cf",x"4a",x"73",x"81"),
  1787 => (x"c3",x"92",x"c2",x"9a"),
  1788 => (x"70",x"30",x"72",x"48"),
  1789 => (x"b0",x"69",x"48",x"4a"),
  1790 => (x"f0",x"c1",x"79",x"70"),
  1791 => (x"78",x"c0",x"48",x"e6"),
  1792 => (x"48",x"e2",x"f0",x"c1"),
  1793 => (x"f6",x"c2",x"78",x"c0"),
  1794 => (x"e4",x"f9",x"49",x"d2"),
  1795 => (x"c0",x"4a",x"70",x"87"),
  1796 => (x"fd",x"03",x"aa",x"b7"),
  1797 => (x"48",x"c0",x"87",x"de"),
  1798 => (x"4d",x"26",x"87",x"c2"),
  1799 => (x"4b",x"26",x"4c",x"26"),
  1800 => (x"00",x"00",x"4f",x"26"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"71",x"1e",x"00",x"00"),
  1803 => (x"ec",x"fc",x"49",x"4a"),
  1804 => (x"1e",x"4f",x"26",x"87"),
  1805 => (x"49",x"72",x"4a",x"c0"),
  1806 => (x"f2",x"c1",x"91",x"c4"),
  1807 => (x"79",x"c0",x"81",x"c2"),
  1808 => (x"b7",x"d0",x"82",x"c1"),
  1809 => (x"87",x"ee",x"04",x"aa"),
  1810 => (x"5e",x"0e",x"4f",x"26"),
  1811 => (x"0e",x"5d",x"5c",x"5b"),
  1812 => (x"cc",x"f8",x"4d",x"71"),
  1813 => (x"c4",x"4a",x"75",x"87"),
  1814 => (x"c1",x"92",x"2a",x"b7"),
  1815 => (x"75",x"82",x"c2",x"f2"),
  1816 => (x"c2",x"9c",x"cf",x"4c"),
  1817 => (x"4b",x"49",x"6a",x"94"),
  1818 => (x"9b",x"c3",x"2b",x"74"),
  1819 => (x"30",x"74",x"48",x"c2"),
  1820 => (x"bc",x"ff",x"4c",x"70"),
  1821 => (x"98",x"71",x"48",x"74"),
  1822 => (x"dc",x"f7",x"7a",x"70"),
  1823 => (x"fe",x"48",x"73",x"87"),
  1824 => (x"00",x"00",x"87",x"d8"),
  1825 => (x"00",x"00",x"00",x"00"),
  1826 => (x"00",x"00",x"00",x"00"),
  1827 => (x"00",x"00",x"00",x"00"),
  1828 => (x"00",x"00",x"00",x"00"),
  1829 => (x"00",x"00",x"00",x"00"),
  1830 => (x"00",x"00",x"00",x"00"),
  1831 => (x"00",x"00",x"00",x"00"),
  1832 => (x"00",x"00",x"00",x"00"),
  1833 => (x"00",x"00",x"00",x"00"),
  1834 => (x"00",x"00",x"00",x"00"),
  1835 => (x"00",x"00",x"00",x"00"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"00",x"00",x"00",x"00"),
  1838 => (x"00",x"00",x"00",x"00"),
  1839 => (x"00",x"00",x"00",x"00"),
  1840 => (x"ff",x"1e",x"00",x"00"),
  1841 => (x"e1",x"c8",x"48",x"d0"),
  1842 => (x"ff",x"48",x"71",x"78"),
  1843 => (x"c4",x"78",x"08",x"d4"),
  1844 => (x"d4",x"ff",x"48",x"66"),
  1845 => (x"4f",x"26",x"78",x"08"),
  1846 => (x"c4",x"4a",x"71",x"1e"),
  1847 => (x"72",x"1e",x"49",x"66"),
  1848 => (x"87",x"de",x"ff",x"49"),
  1849 => (x"c0",x"48",x"d0",x"ff"),
  1850 => (x"26",x"26",x"78",x"e0"),
  1851 => (x"1e",x"73",x"1e",x"4f"),
  1852 => (x"66",x"c8",x"4b",x"71"),
  1853 => (x"4a",x"73",x"1e",x"49"),
  1854 => (x"49",x"a2",x"e0",x"c1"),
  1855 => (x"26",x"87",x"d9",x"ff"),
  1856 => (x"4d",x"26",x"87",x"c4"),
  1857 => (x"4b",x"26",x"4c",x"26"),
  1858 => (x"ff",x"1e",x"4f",x"26"),
  1859 => (x"ff",x"c3",x"4a",x"d4"),
  1860 => (x"48",x"d0",x"ff",x"7a"),
  1861 => (x"de",x"78",x"e1",x"c0"),
  1862 => (x"dc",x"f6",x"c2",x"7a"),
  1863 => (x"48",x"49",x"7a",x"bf"),
  1864 => (x"7a",x"70",x"28",x"c8"),
  1865 => (x"28",x"d0",x"48",x"71"),
  1866 => (x"48",x"71",x"7a",x"70"),
  1867 => (x"7a",x"70",x"28",x"d8"),
  1868 => (x"c0",x"48",x"d0",x"ff"),
  1869 => (x"4f",x"26",x"78",x"e0"),
  1870 => (x"5c",x"5b",x"5e",x"0e"),
  1871 => (x"4c",x"71",x"0e",x"5d"),
  1872 => (x"bf",x"dc",x"f6",x"c2"),
  1873 => (x"2b",x"74",x"4b",x"4d"),
  1874 => (x"c1",x"9b",x"66",x"d0"),
  1875 => (x"ab",x"66",x"d4",x"83"),
  1876 => (x"c0",x"87",x"c2",x"04"),
  1877 => (x"d0",x"4a",x"74",x"4b"),
  1878 => (x"31",x"72",x"49",x"66"),
  1879 => (x"99",x"75",x"b9",x"ff"),
  1880 => (x"30",x"72",x"48",x"73"),
  1881 => (x"71",x"48",x"4a",x"70"),
  1882 => (x"e0",x"f6",x"c2",x"b0"),
  1883 => (x"87",x"da",x"fe",x"58"),
  1884 => (x"4c",x"26",x"4d",x"26"),
  1885 => (x"4f",x"26",x"4b",x"26"),
  1886 => (x"5c",x"5b",x"5e",x"0e"),
  1887 => (x"71",x"1e",x"0e",x"5d"),
  1888 => (x"e0",x"f6",x"c2",x"4c"),
  1889 => (x"c0",x"4a",x"c0",x"4b"),
  1890 => (x"cc",x"fe",x"49",x"f4"),
  1891 => (x"1e",x"74",x"87",x"ea"),
  1892 => (x"49",x"e0",x"f6",x"c2"),
  1893 => (x"87",x"ed",x"e7",x"fe"),
  1894 => (x"49",x"70",x"86",x"c4"),
  1895 => (x"ea",x"c0",x"02",x"99"),
  1896 => (x"a6",x"1e",x"c4",x"87"),
  1897 => (x"f6",x"c2",x"1e",x"4d"),
  1898 => (x"ef",x"fe",x"49",x"e0"),
  1899 => (x"86",x"c8",x"87",x"c4"),
  1900 => (x"d6",x"02",x"98",x"70"),
  1901 => (x"c1",x"4a",x"75",x"87"),
  1902 => (x"c4",x"49",x"c1",x"f8"),
  1903 => (x"e9",x"ca",x"fe",x"4b"),
  1904 => (x"02",x"98",x"70",x"87"),
  1905 => (x"48",x"c0",x"87",x"ca"),
  1906 => (x"c0",x"87",x"ed",x"c0"),
  1907 => (x"87",x"e8",x"c0",x"48"),
  1908 => (x"c1",x"87",x"f3",x"c0"),
  1909 => (x"98",x"70",x"87",x"c4"),
  1910 => (x"c0",x"87",x"c8",x"02"),
  1911 => (x"98",x"70",x"87",x"fc"),
  1912 => (x"c2",x"87",x"f8",x"05"),
  1913 => (x"02",x"bf",x"c0",x"f7"),
  1914 => (x"f6",x"c2",x"87",x"cc"),
  1915 => (x"f7",x"c2",x"48",x"dc"),
  1916 => (x"fc",x"78",x"bf",x"c0"),
  1917 => (x"48",x"c1",x"87",x"d4"),
  1918 => (x"26",x"4d",x"26",x"26"),
  1919 => (x"26",x"4b",x"26",x"4c"),
  1920 => (x"52",x"41",x"5b",x"4f"),
  1921 => (x"c0",x"1e",x"00",x"43"),
  1922 => (x"e0",x"f6",x"c2",x"1e"),
  1923 => (x"f6",x"eb",x"fe",x"49"),
  1924 => (x"f8",x"f6",x"c2",x"87"),
  1925 => (x"26",x"78",x"c0",x"48"),
  1926 => (x"5e",x"0e",x"4f",x"26"),
  1927 => (x"0e",x"5d",x"5c",x"5b"),
  1928 => (x"7e",x"c0",x"86",x"f4"),
  1929 => (x"bf",x"f8",x"f6",x"c2"),
  1930 => (x"a8",x"b7",x"c3",x"48"),
  1931 => (x"c2",x"87",x"d1",x"03"),
  1932 => (x"48",x"bf",x"f8",x"f6"),
  1933 => (x"f6",x"c2",x"80",x"c1"),
  1934 => (x"fb",x"c0",x"58",x"fc"),
  1935 => (x"87",x"d9",x"c6",x"48"),
  1936 => (x"49",x"e0",x"f6",x"c2"),
  1937 => (x"87",x"fe",x"f0",x"fe"),
  1938 => (x"b7",x"c0",x"4c",x"70"),
  1939 => (x"87",x"c4",x"03",x"ac"),
  1940 => (x"87",x"c5",x"c6",x"48"),
  1941 => (x"bf",x"f8",x"f6",x"c2"),
  1942 => (x"02",x"8a",x"c3",x"4a"),
  1943 => (x"8a",x"c1",x"87",x"d8"),
  1944 => (x"87",x"c7",x"c5",x"02"),
  1945 => (x"f2",x"c2",x"02",x"8a"),
  1946 => (x"c1",x"02",x"8a",x"87"),
  1947 => (x"02",x"8a",x"87",x"cf"),
  1948 => (x"c5",x"87",x"de",x"c3"),
  1949 => (x"4d",x"c0",x"87",x"d9"),
  1950 => (x"75",x"5c",x"a6",x"c8"),
  1951 => (x"c1",x"92",x"c4",x"4a"),
  1952 => (x"c2",x"82",x"f7",x"ff"),
  1953 => (x"75",x"4c",x"f4",x"f6"),
  1954 => (x"4b",x"6c",x"97",x"84"),
  1955 => (x"a3",x"c1",x"4b",x"49"),
  1956 => (x"81",x"6a",x"7c",x"97"),
  1957 => (x"a6",x"cc",x"48",x"11"),
  1958 => (x"48",x"66",x"c4",x"58"),
  1959 => (x"02",x"a8",x"66",x"c8"),
  1960 => (x"97",x"c0",x"87",x"c3"),
  1961 => (x"05",x"66",x"c8",x"7c"),
  1962 => (x"f6",x"c2",x"87",x"c7"),
  1963 => (x"a5",x"c4",x"48",x"f8"),
  1964 => (x"c4",x"85",x"c1",x"78"),
  1965 => (x"ff",x"04",x"ad",x"b7"),
  1966 => (x"d2",x"c4",x"87",x"c1"),
  1967 => (x"c4",x"f7",x"c2",x"87"),
  1968 => (x"b7",x"c8",x"48",x"bf"),
  1969 => (x"87",x"cb",x"01",x"a8"),
  1970 => (x"c6",x"02",x"ac",x"ca"),
  1971 => (x"05",x"ac",x"cd",x"87"),
  1972 => (x"c2",x"87",x"f3",x"c0"),
  1973 => (x"4b",x"bf",x"c4",x"f7"),
  1974 => (x"03",x"ab",x"b7",x"c8"),
  1975 => (x"f7",x"c2",x"87",x"d2"),
  1976 => (x"81",x"73",x"49",x"c8"),
  1977 => (x"c1",x"51",x"e0",x"c0"),
  1978 => (x"ab",x"b7",x"c8",x"83"),
  1979 => (x"87",x"ee",x"ff",x"04"),
  1980 => (x"48",x"d0",x"f7",x"c2"),
  1981 => (x"c1",x"50",x"d2",x"c1"),
  1982 => (x"cd",x"c1",x"50",x"cf"),
  1983 => (x"e4",x"50",x"c0",x"50"),
  1984 => (x"c3",x"78",x"c3",x"80"),
  1985 => (x"f7",x"c2",x"87",x"c9"),
  1986 => (x"48",x"49",x"bf",x"c4"),
  1987 => (x"f7",x"c2",x"80",x"c1"),
  1988 => (x"c4",x"48",x"58",x"c8"),
  1989 => (x"51",x"74",x"81",x"a0"),
  1990 => (x"c0",x"87",x"f4",x"c2"),
  1991 => (x"04",x"ac",x"b7",x"f0"),
  1992 => (x"f9",x"c0",x"87",x"da"),
  1993 => (x"d3",x"01",x"ac",x"b7"),
  1994 => (x"fc",x"f6",x"c2",x"87"),
  1995 => (x"91",x"ca",x"49",x"bf"),
  1996 => (x"f0",x"c0",x"4a",x"74"),
  1997 => (x"fc",x"f6",x"c2",x"8a"),
  1998 => (x"78",x"a1",x"72",x"48"),
  1999 => (x"c0",x"02",x"ac",x"ca"),
  2000 => (x"ac",x"cd",x"87",x"c6"),
  2001 => (x"87",x"c7",x"c2",x"05"),
  2002 => (x"48",x"f8",x"f6",x"c2"),
  2003 => (x"fe",x"c1",x"78",x"c3"),
  2004 => (x"b7",x"f0",x"c0",x"87"),
  2005 => (x"87",x"db",x"04",x"ac"),
  2006 => (x"ac",x"b7",x"f9",x"c0"),
  2007 => (x"87",x"d3",x"c0",x"01"),
  2008 => (x"bf",x"c0",x"f7",x"c2"),
  2009 => (x"74",x"91",x"d0",x"49"),
  2010 => (x"8a",x"f0",x"c0",x"4a"),
  2011 => (x"48",x"c0",x"f7",x"c2"),
  2012 => (x"c1",x"78",x"a1",x"72"),
  2013 => (x"04",x"ac",x"b7",x"c1"),
  2014 => (x"c1",x"87",x"db",x"c0"),
  2015 => (x"01",x"ac",x"b7",x"c6"),
  2016 => (x"c2",x"87",x"d3",x"c0"),
  2017 => (x"49",x"bf",x"c0",x"f7"),
  2018 => (x"4a",x"74",x"91",x"d0"),
  2019 => (x"c2",x"8a",x"f7",x"c0"),
  2020 => (x"72",x"48",x"c0",x"f7"),
  2021 => (x"ac",x"ca",x"78",x"a1"),
  2022 => (x"87",x"c6",x"c0",x"02"),
  2023 => (x"c0",x"05",x"ac",x"cd"),
  2024 => (x"f6",x"c2",x"87",x"ed"),
  2025 => (x"78",x"c3",x"48",x"f8"),
  2026 => (x"c0",x"87",x"e4",x"c0"),
  2027 => (x"c0",x"05",x"ac",x"e2"),
  2028 => (x"fb",x"c0",x"87",x"c6"),
  2029 => (x"87",x"d7",x"c0",x"7e"),
  2030 => (x"c0",x"02",x"ac",x"ca"),
  2031 => (x"ac",x"cd",x"87",x"c6"),
  2032 => (x"87",x"c9",x"c0",x"05"),
  2033 => (x"48",x"f8",x"f6",x"c2"),
  2034 => (x"c2",x"c0",x"78",x"c3"),
  2035 => (x"6e",x"7e",x"74",x"87"),
  2036 => (x"87",x"d0",x"f9",x"02"),
  2037 => (x"ff",x"c3",x"48",x"6e"),
  2038 => (x"f8",x"8e",x"f4",x"99"),
  2039 => (x"4f",x"43",x"87",x"db"),
  2040 => (x"00",x"3d",x"46",x"4e"),
  2041 => (x"00",x"44",x"4f",x"4d"),
  2042 => (x"45",x"4d",x"41",x"4e"),
  2043 => (x"46",x"45",x"44",x"00"),
  2044 => (x"54",x"4c",x"55",x"41"),
  2045 => (x"de",x"00",x"30",x"3d"),
  2046 => (x"e4",x"00",x"00",x"1f"),
  2047 => (x"e8",x"00",x"00",x"1f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

