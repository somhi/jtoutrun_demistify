library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"00444f4d",
     1 => x"454d414e",
     2 => x"46454400",
     3 => x"544c5541",
     4 => x"fa00303d",
     5 => x"0000001f",
     6 => x"04000020",
     7 => x"09000020",
     8 => x"1e000020",
     9 => x"c848d0ff",
    10 => x"487178c9",
    11 => x"7808d4ff",
    12 => x"711e4f26",
    13 => x"87eb494a",
    14 => x"c848d0ff",
    15 => x"1e4f2678",
    16 => x"4b711e73",
    17 => x"bff8f9c2",
    18 => x"c287c302",
    19 => x"d0ff87eb",
    20 => x"78c9c848",
    21 => x"e0c04973",
    22 => x"48d4ffb1",
    23 => x"f9c27871",
    24 => x"78c048ec",
    25 => x"c50266c8",
    26 => x"49ffc387",
    27 => x"49c087c2",
    28 => x"59f4f9c2",
    29 => x"c60266cc",
    30 => x"d5d5c587",
    31 => x"cf87c44a",
    32 => x"c24affff",
    33 => x"c25af8f9",
    34 => x"c148f8f9",
    35 => x"2687c478",
    36 => x"264c264d",
    37 => x"0e4f264b",
    38 => x"5d5c5b5e",
    39 => x"c24a710e",
    40 => x"4cbff4f9",
    41 => x"cb029a72",
    42 => x"91c84987",
    43 => x"4bf5c0c2",
    44 => x"87c48371",
    45 => x"4bf5c4c2",
    46 => x"49134dc0",
    47 => x"f9c29974",
    48 => x"ffb9bff0",
    49 => x"787148d4",
    50 => x"852cb7c1",
    51 => x"04adb7c8",
    52 => x"f9c287e8",
    53 => x"c848bfec",
    54 => x"f0f9c280",
    55 => x"87effe58",
    56 => x"711e731e",
    57 => x"9a4a134b",
    58 => x"7287cb02",
    59 => x"87e7fe49",
    60 => x"059a4a13",
    61 => x"dafe87f5",
    62 => x"f9c21e87",
    63 => x"c249bfec",
    64 => x"c148ecf9",
    65 => x"c0c478a1",
    66 => x"db03a9b7",
    67 => x"48d4ff87",
    68 => x"bff0f9c2",
    69 => x"ecf9c278",
    70 => x"f9c249bf",
    71 => x"a1c148ec",
    72 => x"b7c0c478",
    73 => x"87e504a9",
    74 => x"c848d0ff",
    75 => x"f8f9c278",
    76 => x"2678c048",
    77 => x"0000004f",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"00005f5f",
    81 => x"03030000",
    82 => x"00030300",
    83 => x"7f7f1400",
    84 => x"147f7f14",
    85 => x"2e240000",
    86 => x"123a6b6b",
    87 => x"366a4c00",
    88 => x"32566c18",
    89 => x"4f7e3000",
    90 => x"683a7759",
    91 => x"04000040",
    92 => x"00000307",
    93 => x"1c000000",
    94 => x"0041633e",
    95 => x"41000000",
    96 => x"001c3e63",
    97 => x"3e2a0800",
    98 => x"2a3e1c1c",
    99 => x"08080008",
   100 => x"08083e3e",
   101 => x"80000000",
   102 => x"000060e0",
   103 => x"08080000",
   104 => x"08080808",
   105 => x"00000000",
   106 => x"00006060",
   107 => x"30604000",
   108 => x"03060c18",
   109 => x"7f3e0001",
   110 => x"3e7f4d59",
   111 => x"06040000",
   112 => x"00007f7f",
   113 => x"63420000",
   114 => x"464f5971",
   115 => x"63220000",
   116 => x"367f4949",
   117 => x"161c1800",
   118 => x"107f7f13",
   119 => x"67270000",
   120 => x"397d4545",
   121 => x"7e3c0000",
   122 => x"3079494b",
   123 => x"01010000",
   124 => x"070f7971",
   125 => x"7f360000",
   126 => x"367f4949",
   127 => x"4f060000",
   128 => x"1e3f6949",
   129 => x"00000000",
   130 => x"00006666",
   131 => x"80000000",
   132 => x"000066e6",
   133 => x"08080000",
   134 => x"22221414",
   135 => x"14140000",
   136 => x"14141414",
   137 => x"22220000",
   138 => x"08081414",
   139 => x"03020000",
   140 => x"060f5951",
   141 => x"417f3e00",
   142 => x"1e1f555d",
   143 => x"7f7e0000",
   144 => x"7e7f0909",
   145 => x"7f7f0000",
   146 => x"367f4949",
   147 => x"3e1c0000",
   148 => x"41414163",
   149 => x"7f7f0000",
   150 => x"1c3e6341",
   151 => x"7f7f0000",
   152 => x"41414949",
   153 => x"7f7f0000",
   154 => x"01010909",
   155 => x"7f3e0000",
   156 => x"7a7b4941",
   157 => x"7f7f0000",
   158 => x"7f7f0808",
   159 => x"41000000",
   160 => x"00417f7f",
   161 => x"60200000",
   162 => x"3f7f4040",
   163 => x"087f7f00",
   164 => x"4163361c",
   165 => x"7f7f0000",
   166 => x"40404040",
   167 => x"067f7f00",
   168 => x"7f7f060c",
   169 => x"067f7f00",
   170 => x"7f7f180c",
   171 => x"7f3e0000",
   172 => x"3e7f4141",
   173 => x"7f7f0000",
   174 => x"060f0909",
   175 => x"417f3e00",
   176 => x"407e7f61",
   177 => x"7f7f0000",
   178 => x"667f1909",
   179 => x"6f260000",
   180 => x"327b594d",
   181 => x"01010000",
   182 => x"01017f7f",
   183 => x"7f3f0000",
   184 => x"3f7f4040",
   185 => x"3f0f0000",
   186 => x"0f3f7070",
   187 => x"307f7f00",
   188 => x"7f7f3018",
   189 => x"36634100",
   190 => x"63361c1c",
   191 => x"06030141",
   192 => x"03067c7c",
   193 => x"59716101",
   194 => x"4143474d",
   195 => x"7f000000",
   196 => x"0041417f",
   197 => x"06030100",
   198 => x"6030180c",
   199 => x"41000040",
   200 => x"007f7f41",
   201 => x"060c0800",
   202 => x"080c0603",
   203 => x"80808000",
   204 => x"80808080",
   205 => x"00000000",
   206 => x"00040703",
   207 => x"74200000",
   208 => x"787c5454",
   209 => x"7f7f0000",
   210 => x"387c4444",
   211 => x"7c380000",
   212 => x"00444444",
   213 => x"7c380000",
   214 => x"7f7f4444",
   215 => x"7c380000",
   216 => x"185c5454",
   217 => x"7e040000",
   218 => x"0005057f",
   219 => x"bc180000",
   220 => x"7cfca4a4",
   221 => x"7f7f0000",
   222 => x"787c0404",
   223 => x"00000000",
   224 => x"00407d3d",
   225 => x"80800000",
   226 => x"007dfd80",
   227 => x"7f7f0000",
   228 => x"446c3810",
   229 => x"00000000",
   230 => x"00407f3f",
   231 => x"0c7c7c00",
   232 => x"787c0c18",
   233 => x"7c7c0000",
   234 => x"787c0404",
   235 => x"7c380000",
   236 => x"387c4444",
   237 => x"fcfc0000",
   238 => x"183c2424",
   239 => x"3c180000",
   240 => x"fcfc2424",
   241 => x"7c7c0000",
   242 => x"080c0404",
   243 => x"5c480000",
   244 => x"20745454",
   245 => x"3f040000",
   246 => x"0044447f",
   247 => x"7c3c0000",
   248 => x"7c7c4040",
   249 => x"3c1c0000",
   250 => x"1c3c6060",
   251 => x"607c3c00",
   252 => x"3c7c6030",
   253 => x"386c4400",
   254 => x"446c3810",
   255 => x"bc1c0000",
   256 => x"1c3c60e0",
   257 => x"64440000",
   258 => x"444c5c74",
   259 => x"08080000",
   260 => x"4141773e",
   261 => x"00000000",
   262 => x"00007f7f",
   263 => x"41410000",
   264 => x"08083e77",
   265 => x"01010200",
   266 => x"01020203",
   267 => x"7f7f7f00",
   268 => x"7f7f7f7f",
   269 => x"1c080800",
   270 => x"7f3e3e1c",
   271 => x"3e7f7f7f",
   272 => x"081c1c3e",
   273 => x"18100008",
   274 => x"10187c7c",
   275 => x"30100000",
   276 => x"10307c7c",
   277 => x"60301000",
   278 => x"061e7860",
   279 => x"3c664200",
   280 => x"42663c18",
   281 => x"6a387800",
   282 => x"386cc6c2",
   283 => x"00006000",
   284 => x"60000060",
   285 => x"5b5e0e00",
   286 => x"1e0e5d5c",
   287 => x"fac24c71",
   288 => x"c04dbfc9",
   289 => x"741ec04b",
   290 => x"87c702ab",
   291 => x"c048a6c4",
   292 => x"c487c578",
   293 => x"78c148a6",
   294 => x"731e66c4",
   295 => x"87dfee49",
   296 => x"e0c086c8",
   297 => x"87efef49",
   298 => x"6a4aa5c4",
   299 => x"87f0f049",
   300 => x"cb87c6f1",
   301 => x"c883c185",
   302 => x"ff04abb7",
   303 => x"262687c7",
   304 => x"264c264d",
   305 => x"1e4f264b",
   306 => x"fac24a71",
   307 => x"fac25acd",
   308 => x"78c748cd",
   309 => x"87ddfe49",
   310 => x"731e4f26",
   311 => x"c04a711e",
   312 => x"d303aab7",
   313 => x"fae0c287",
   314 => x"87c405bf",
   315 => x"87c24bc1",
   316 => x"e0c24bc0",
   317 => x"87c45bfe",
   318 => x"5afee0c2",
   319 => x"bffae0c2",
   320 => x"c19ac14a",
   321 => x"ec49a2c0",
   322 => x"48fc87e8",
   323 => x"bffae0c2",
   324 => x"87effe78",
   325 => x"c44a711e",
   326 => x"49721e66",
   327 => x"87dddfff",
   328 => x"1e4f2626",
   329 => x"bffae0c2",
   330 => x"cddcff49",
   331 => x"c1fac287",
   332 => x"78bfe848",
   333 => x"48fdf9c2",
   334 => x"c278bfec",
   335 => x"4abfc1fa",
   336 => x"99ffc349",
   337 => x"722ab7c8",
   338 => x"c2b07148",
   339 => x"2658c9fa",
   340 => x"5b5e0e4f",
   341 => x"710e5d5c",
   342 => x"87c7ff4b",
   343 => x"48fcf9c2",
   344 => x"497350c0",
   345 => x"87f2dbff",
   346 => x"c24c4970",
   347 => x"49eecb9c",
   348 => x"7087cfcb",
   349 => x"f9c24d49",
   350 => x"05bf97fc",
   351 => x"d087e4c1",
   352 => x"fac24966",
   353 => x"0599bfc5",
   354 => x"66d487d7",
   355 => x"fdf9c249",
   356 => x"cc0599bf",
   357 => x"ff497387",
   358 => x"7087ffda",
   359 => x"c2c10298",
   360 => x"fd4cc187",
   361 => x"497587fd",
   362 => x"7087e3ca",
   363 => x"87c60298",
   364 => x"48fcf9c2",
   365 => x"f9c250c1",
   366 => x"05bf97fc",
   367 => x"c287e4c0",
   368 => x"49bfc5fa",
   369 => x"059966d0",
   370 => x"c287d6ff",
   371 => x"49bffdf9",
   372 => x"059966d4",
   373 => x"7387caff",
   374 => x"fdd9ff49",
   375 => x"05987087",
   376 => x"7487fefe",
   377 => x"87d7fb48",
   378 => x"5c5b5e0e",
   379 => x"86f40e5d",
   380 => x"ec4c4dc0",
   381 => x"a6c47ebf",
   382 => x"c9fac248",
   383 => x"1ec178bf",
   384 => x"49c71ec0",
   385 => x"c887cafd",
   386 => x"02987086",
   387 => x"49ff87ce",
   388 => x"c187c7fb",
   389 => x"d9ff49da",
   390 => x"4dc187c0",
   391 => x"97fcf9c2",
   392 => x"87c302bf",
   393 => x"c287c0c9",
   394 => x"4bbfc1fa",
   395 => x"bffae0c2",
   396 => x"87ebc005",
   397 => x"ff49fdc3",
   398 => x"c387dfd8",
   399 => x"d8ff49fa",
   400 => x"497387d8",
   401 => x"7199ffc3",
   402 => x"fb49c01e",
   403 => x"497387c6",
   404 => x"7129b7c8",
   405 => x"fa49c11e",
   406 => x"86c887fa",
   407 => x"c287c1c6",
   408 => x"4bbfc5fa",
   409 => x"87dd029b",
   410 => x"bff6e0c2",
   411 => x"87dec749",
   412 => x"c4059870",
   413 => x"d24bc087",
   414 => x"49e0c287",
   415 => x"c287c3c7",
   416 => x"c658fae0",
   417 => x"f6e0c287",
   418 => x"7378c048",
   419 => x"0599c249",
   420 => x"ebc387ce",
   421 => x"c1d7ff49",
   422 => x"c2497087",
   423 => x"87c20299",
   424 => x"49734cfb",
   425 => x"ce0599c1",
   426 => x"49f4c387",
   427 => x"87ead6ff",
   428 => x"99c24970",
   429 => x"fa87c202",
   430 => x"c849734c",
   431 => x"87ce0599",
   432 => x"ff49f5c3",
   433 => x"7087d3d6",
   434 => x"0299c249",
   435 => x"fac287d5",
   436 => x"ca02bfcd",
   437 => x"88c14887",
   438 => x"58d1fac2",
   439 => x"ff87c2c0",
   440 => x"734dc14c",
   441 => x"0599c449",
   442 => x"f2c387ce",
   443 => x"e9d5ff49",
   444 => x"c2497087",
   445 => x"87dc0299",
   446 => x"bfcdfac2",
   447 => x"b7c7487e",
   448 => x"cbc003a8",
   449 => x"c1486e87",
   450 => x"d1fac280",
   451 => x"87c2c058",
   452 => x"4dc14cfe",
   453 => x"ff49fdc3",
   454 => x"7087ffd4",
   455 => x"0299c249",
   456 => x"c287d5c0",
   457 => x"02bfcdfa",
   458 => x"c287c9c0",
   459 => x"c048cdfa",
   460 => x"87c2c078",
   461 => x"4dc14cfd",
   462 => x"ff49fac3",
   463 => x"7087dbd4",
   464 => x"0299c249",
   465 => x"c287d9c0",
   466 => x"48bfcdfa",
   467 => x"03a8b7c7",
   468 => x"c287c9c0",
   469 => x"c748cdfa",
   470 => x"87c2c078",
   471 => x"4dc14cfc",
   472 => x"03acb7c0",
   473 => x"c487d1c0",
   474 => x"d8c14a66",
   475 => x"c0026a82",
   476 => x"4b6a87c6",
   477 => x"0f734974",
   478 => x"f0c31ec0",
   479 => x"49dac11e",
   480 => x"c887cef7",
   481 => x"02987086",
   482 => x"c887e2c0",
   483 => x"fac248a6",
   484 => x"c878bfcd",
   485 => x"91cb4966",
   486 => x"714866c4",
   487 => x"6e7e7080",
   488 => x"c8c002bf",
   489 => x"4bbf6e87",
   490 => x"734966c8",
   491 => x"029d750f",
   492 => x"c287c8c0",
   493 => x"49bfcdfa",
   494 => x"c287faf2",
   495 => x"02bffee0",
   496 => x"4987ddc0",
   497 => x"7087c7c2",
   498 => x"d3c00298",
   499 => x"cdfac287",
   500 => x"e0f249bf",
   501 => x"f449c087",
   502 => x"e0c287c0",
   503 => x"78c048fe",
   504 => x"daf38ef4",
   505 => x"5b5e0e87",
   506 => x"1e0e5d5c",
   507 => x"fac24c71",
   508 => x"c149bfc9",
   509 => x"c14da1cd",
   510 => x"7e6981d1",
   511 => x"cf029c74",
   512 => x"4ba5c487",
   513 => x"fac27b74",
   514 => x"f249bfc9",
   515 => x"7b6e87f9",
   516 => x"c4059c74",
   517 => x"c24bc087",
   518 => x"734bc187",
   519 => x"87faf249",
   520 => x"c70266d4",
   521 => x"87da4987",
   522 => x"87c24a70",
   523 => x"e1c24ac0",
   524 => x"f2265ac2",
   525 => x"000087c9",
   526 => x"00000000",
   527 => x"00000000",
   528 => x"711e0000",
   529 => x"bfc8ff4a",
   530 => x"48a17249",
   531 => x"ff1e4f26",
   532 => x"fe89bfc8",
   533 => x"c0c0c0c0",
   534 => x"c401a9c0",
   535 => x"c24ac087",
   536 => x"724ac187",
   537 => x"1e4f2648",
   538 => x"bff5e2c2",
   539 => x"c2b9c149",
   540 => x"ff59f9e2",
   541 => x"ffc348d4",
   542 => x"48d0ff78",
   543 => x"ff78e1c0",
   544 => x"78c148d4",
   545 => x"787131c4",
   546 => x"c048d0ff",
   547 => x"4f2678e0",
   548 => x"e9e2c21e",
   549 => x"f0f4c21e",
   550 => x"d4fdfd49",
   551 => x"7086c487",
   552 => x"87c30298",
   553 => x"2687c0ff",
   554 => x"4b35314f",
   555 => x"20205a48",
   556 => x"47464320",
   557 => x"00000000",
   558 => x"5b5e0e00",
   559 => x"c20e5d5c",
   560 => x"4abffdf9",
   561 => x"bfe2e4c2",
   562 => x"bc724c49",
   563 => x"c6ff4d71",
   564 => x"4bc087de",
   565 => x"99d04974",
   566 => x"87e7c002",
   567 => x"c848d0ff",
   568 => x"d4ff78e1",
   569 => x"7578c548",
   570 => x"0299d049",
   571 => x"f0c387c3",
   572 => x"cae7c278",
   573 => x"11817349",
   574 => x"08d4ff48",
   575 => x"48d0ff78",
   576 => x"c178e0c0",
   577 => x"c8832d2c",
   578 => x"c7ff04ab",
   579 => x"d7c5ff87",
   580 => x"e2e4c287",
   581 => x"fdf9c248",
   582 => x"4d2678bf",
   583 => x"4b264c26",
   584 => x"00004f26",
   585 => x"731e0000",
   586 => x"c14bc01e",
   587 => x"de48d7e7",
   588 => x"c21ec850",
   589 => x"fe49d1fa",
   590 => x"c487c1d5",
   591 => x"c21e7286",
   592 => x"c248d8e6",
   593 => x"c449d9fa",
   594 => x"41204aa1",
   595 => x"f905aa71",
   596 => x"c24a2687",
   597 => x"fd49dce6",
   598 => x"7087f7f8",
   599 => x"c5029a4a",
   600 => x"c7fe4987",
   601 => x"1e7287e0",
   602 => x"48e8e6c2",
   603 => x"49d9fac2",
   604 => x"204aa1c4",
   605 => x"05aa7141",
   606 => x"4a2687f9",
   607 => x"49d1fac2",
   608 => x"87d1d9fe",
   609 => x"c4059870",
   610 => x"ece6c287",
   611 => x"fe49c04b",
   612 => x"7387d5c5",
   613 => x"87c6fe48",
   614 => x"00202020",
   615 => x"45544f4a",
   616 => x"20204f47",
   617 => x"00202020",
   618 => x"00435241",
   619 => x"20435241",
   620 => x"64616f6c",
   621 => x"20676e69",
   622 => x"6c696166",
   623 => x"1e006465",
   624 => x"fb87e5f0",
   625 => x"87f887f3",
   626 => x"1e164f26",
   627 => x"362e2526",
   628 => x"362e3e3d",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
