library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fcf8c287",
    12 => x"86c0c54e",
    13 => x"49fcf8c2",
    14 => x"48fce5c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087ede5",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"711e4f26",
    53 => x"4966c44a",
    54 => x"c888c148",
    55 => x"997158a6",
    56 => x"ff87d602",
    57 => x"ffc348d4",
    58 => x"c4526878",
    59 => x"c1484966",
    60 => x"58a6c888",
    61 => x"ea059971",
    62 => x"1e4f2687",
    63 => x"d4ff1e73",
    64 => x"7bffc34b",
    65 => x"ffc34a6b",
    66 => x"c8496b7b",
    67 => x"c3b17232",
    68 => x"4a6b7bff",
    69 => x"b27131c8",
    70 => x"6b7bffc3",
    71 => x"7232c849",
    72 => x"c44871b1",
    73 => x"264d2687",
    74 => x"264b264c",
    75 => x"5b5e0e4f",
    76 => x"710e5d5c",
    77 => x"4cd4ff4a",
    78 => x"ffc34972",
    79 => x"c27c7199",
    80 => x"05bffce5",
    81 => x"66d087c8",
    82 => x"d430c948",
    83 => x"66d058a6",
    84 => x"c329d849",
    85 => x"7c7199ff",
    86 => x"d04966d0",
    87 => x"99ffc329",
    88 => x"66d07c71",
    89 => x"c329c849",
    90 => x"7c7199ff",
    91 => x"c34966d0",
    92 => x"7c7199ff",
    93 => x"29d04972",
    94 => x"7199ffc3",
    95 => x"c94b6c7c",
    96 => x"c34dfff0",
    97 => x"d005abff",
    98 => x"7cffc387",
    99 => x"8dc14b6c",
   100 => x"c387c602",
   101 => x"f002abff",
   102 => x"fe487387",
   103 => x"c01e87c7",
   104 => x"48d4ff49",
   105 => x"c178ffc3",
   106 => x"b7c8c381",
   107 => x"87f104a9",
   108 => x"731e4f26",
   109 => x"c487e71e",
   110 => x"c04bdff8",
   111 => x"f0ffc01e",
   112 => x"fd49f7c1",
   113 => x"86c487e7",
   114 => x"c005a8c1",
   115 => x"d4ff87ea",
   116 => x"78ffc348",
   117 => x"c0c0c0c1",
   118 => x"c01ec0c0",
   119 => x"e9c1f0e1",
   120 => x"87c9fd49",
   121 => x"987086c4",
   122 => x"ff87ca05",
   123 => x"ffc348d4",
   124 => x"cb48c178",
   125 => x"87e6fe87",
   126 => x"fe058bc1",
   127 => x"48c087fd",
   128 => x"1e87e6fc",
   129 => x"d4ff1e73",
   130 => x"78ffc348",
   131 => x"1ec04bd3",
   132 => x"c1f0ffc0",
   133 => x"d4fc49c1",
   134 => x"7086c487",
   135 => x"87ca0598",
   136 => x"c348d4ff",
   137 => x"48c178ff",
   138 => x"f1fd87cb",
   139 => x"058bc187",
   140 => x"c087dbff",
   141 => x"87f1fb48",
   142 => x"5c5b5e0e",
   143 => x"4cd4ff0e",
   144 => x"c687dbfd",
   145 => x"e1c01eea",
   146 => x"49c8c1f0",
   147 => x"c487defb",
   148 => x"02a8c186",
   149 => x"eafe87c8",
   150 => x"c148c087",
   151 => x"dafa87e2",
   152 => x"cf497087",
   153 => x"c699ffff",
   154 => x"c802a9ea",
   155 => x"87d3fe87",
   156 => x"cbc148c0",
   157 => x"7cffc387",
   158 => x"fc4bf1c0",
   159 => x"987087f4",
   160 => x"87ebc002",
   161 => x"ffc01ec0",
   162 => x"49fac1f0",
   163 => x"c487defa",
   164 => x"05987086",
   165 => x"ffc387d9",
   166 => x"c3496c7c",
   167 => x"7c7c7cff",
   168 => x"99c0c17c",
   169 => x"c187c402",
   170 => x"c087d548",
   171 => x"c287d148",
   172 => x"87c405ab",
   173 => x"87c848c0",
   174 => x"fe058bc1",
   175 => x"48c087fd",
   176 => x"1e87e4f9",
   177 => x"e5c21e73",
   178 => x"78c148fc",
   179 => x"d0ff4bc7",
   180 => x"fb78c248",
   181 => x"d0ff87c8",
   182 => x"c078c348",
   183 => x"d0e5c01e",
   184 => x"f949c0c1",
   185 => x"86c487c7",
   186 => x"c105a8c1",
   187 => x"abc24b87",
   188 => x"c087c505",
   189 => x"87f9c048",
   190 => x"ff058bc1",
   191 => x"f7fc87d0",
   192 => x"c0e6c287",
   193 => x"05987058",
   194 => x"1ec187cd",
   195 => x"c1f0ffc0",
   196 => x"d8f849d0",
   197 => x"ff86c487",
   198 => x"ffc348d4",
   199 => x"87fcc278",
   200 => x"58c4e6c2",
   201 => x"c248d0ff",
   202 => x"48d4ff78",
   203 => x"c178ffc3",
   204 => x"87f5f748",
   205 => x"5c5b5e0e",
   206 => x"4b710e5d",
   207 => x"eec54cc0",
   208 => x"ff4adfcd",
   209 => x"ffc348d4",
   210 => x"c3496878",
   211 => x"c005a9fe",
   212 => x"4d7087fd",
   213 => x"cc029b73",
   214 => x"1e66d087",
   215 => x"f1f54973",
   216 => x"d686c487",
   217 => x"48d0ff87",
   218 => x"c378d1c4",
   219 => x"66d07dff",
   220 => x"d488c148",
   221 => x"987058a6",
   222 => x"ff87f005",
   223 => x"ffc348d4",
   224 => x"9b737878",
   225 => x"ff87c505",
   226 => x"78d048d0",
   227 => x"c14c4ac1",
   228 => x"eefe058a",
   229 => x"f6487487",
   230 => x"731e87cb",
   231 => x"c04a711e",
   232 => x"48d4ff4b",
   233 => x"ff78ffc3",
   234 => x"c3c448d0",
   235 => x"48d4ff78",
   236 => x"7278ffc3",
   237 => x"f0ffc01e",
   238 => x"f549d1c1",
   239 => x"86c487ef",
   240 => x"d2059870",
   241 => x"1ec0c887",
   242 => x"fd4966cc",
   243 => x"86c487e6",
   244 => x"d0ff4b70",
   245 => x"7378c248",
   246 => x"87cdf548",
   247 => x"5c5b5e0e",
   248 => x"1ec00e5d",
   249 => x"c1f0ffc0",
   250 => x"c0f549c9",
   251 => x"c21ed287",
   252 => x"fc49c4e6",
   253 => x"86c887fe",
   254 => x"84c14cc0",
   255 => x"04acb7d2",
   256 => x"e6c287f8",
   257 => x"49bf97c4",
   258 => x"c199c0c3",
   259 => x"c005a9c0",
   260 => x"e6c287e7",
   261 => x"49bf97cb",
   262 => x"e6c231d0",
   263 => x"4abf97cc",
   264 => x"b17232c8",
   265 => x"97cde6c2",
   266 => x"71b14abf",
   267 => x"ffffcf4c",
   268 => x"84c19cff",
   269 => x"e7c134ca",
   270 => x"cde6c287",
   271 => x"c149bf97",
   272 => x"c299c631",
   273 => x"bf97cee6",
   274 => x"2ab7c74a",
   275 => x"e6c2b172",
   276 => x"4abf97c9",
   277 => x"c29dcf4d",
   278 => x"bf97cae6",
   279 => x"ca9ac34a",
   280 => x"cbe6c232",
   281 => x"c24bbf97",
   282 => x"c2b27333",
   283 => x"bf97cce6",
   284 => x"9bc0c34b",
   285 => x"732bb7c6",
   286 => x"c181c2b2",
   287 => x"70307148",
   288 => x"7548c149",
   289 => x"724d7030",
   290 => x"7184c14c",
   291 => x"b7c0c894",
   292 => x"87cc06ad",
   293 => x"2db734c1",
   294 => x"adb7c0c8",
   295 => x"87f4ff01",
   296 => x"c0f24874",
   297 => x"5b5e0e87",
   298 => x"f80e5d5c",
   299 => x"eaeec286",
   300 => x"c278c048",
   301 => x"c01ee2e6",
   302 => x"87defb49",
   303 => x"987086c4",
   304 => x"c087c505",
   305 => x"87cec948",
   306 => x"7ec14dc0",
   307 => x"bfe1f5c0",
   308 => x"d8e7c249",
   309 => x"4bc8714a",
   310 => x"7087cfee",
   311 => x"87c20598",
   312 => x"f5c07ec0",
   313 => x"c249bfdd",
   314 => x"714af4e7",
   315 => x"f9ed4bc8",
   316 => x"05987087",
   317 => x"7ec087c2",
   318 => x"fdc0026e",
   319 => x"e8edc287",
   320 => x"eec24dbf",
   321 => x"7ebf9fe0",
   322 => x"ead6c548",
   323 => x"87c705a8",
   324 => x"bfe8edc2",
   325 => x"6e87ce4d",
   326 => x"d5e9ca48",
   327 => x"87c502a8",
   328 => x"f1c748c0",
   329 => x"e2e6c287",
   330 => x"f949751e",
   331 => x"86c487ec",
   332 => x"c5059870",
   333 => x"c748c087",
   334 => x"f5c087dc",
   335 => x"c249bfdd",
   336 => x"714af4e7",
   337 => x"e1ec4bc8",
   338 => x"05987087",
   339 => x"eec287c8",
   340 => x"78c148ea",
   341 => x"f5c087da",
   342 => x"c249bfe1",
   343 => x"714ad8e7",
   344 => x"c5ec4bc8",
   345 => x"02987087",
   346 => x"c087c5c0",
   347 => x"87e6c648",
   348 => x"97e0eec2",
   349 => x"d5c149bf",
   350 => x"cdc005a9",
   351 => x"e1eec287",
   352 => x"c249bf97",
   353 => x"c002a9ea",
   354 => x"48c087c5",
   355 => x"c287c7c6",
   356 => x"bf97e2e6",
   357 => x"e9c3487e",
   358 => x"cec002a8",
   359 => x"c3486e87",
   360 => x"c002a8eb",
   361 => x"48c087c5",
   362 => x"c287ebc5",
   363 => x"bf97ede6",
   364 => x"c0059949",
   365 => x"e6c287cc",
   366 => x"49bf97ee",
   367 => x"c002a9c2",
   368 => x"48c087c5",
   369 => x"c287cfc5",
   370 => x"bf97efe6",
   371 => x"e6eec248",
   372 => x"484c7058",
   373 => x"eec288c1",
   374 => x"e6c258ea",
   375 => x"49bf97f0",
   376 => x"e6c28175",
   377 => x"4abf97f1",
   378 => x"a17232c8",
   379 => x"f7f2c27e",
   380 => x"c2786e48",
   381 => x"bf97f2e6",
   382 => x"58a6c848",
   383 => x"bfeaeec2",
   384 => x"87d4c202",
   385 => x"bfddf5c0",
   386 => x"f4e7c249",
   387 => x"4bc8714a",
   388 => x"7087d7e9",
   389 => x"c5c00298",
   390 => x"c348c087",
   391 => x"eec287f8",
   392 => x"c24cbfe2",
   393 => x"c25ccbf3",
   394 => x"bf97c7e7",
   395 => x"c231c849",
   396 => x"bf97c6e7",
   397 => x"c249a14a",
   398 => x"bf97c8e7",
   399 => x"7232d04a",
   400 => x"e7c249a1",
   401 => x"4abf97c9",
   402 => x"a17232d8",
   403 => x"9166c449",
   404 => x"bff7f2c2",
   405 => x"fff2c281",
   406 => x"cfe7c259",
   407 => x"c84abf97",
   408 => x"cee7c232",
   409 => x"a24bbf97",
   410 => x"d0e7c24a",
   411 => x"d04bbf97",
   412 => x"4aa27333",
   413 => x"97d1e7c2",
   414 => x"9bcf4bbf",
   415 => x"a27333d8",
   416 => x"c3f3c24a",
   417 => x"fff2c25a",
   418 => x"8ac24abf",
   419 => x"f3c29274",
   420 => x"a17248c3",
   421 => x"87cac178",
   422 => x"97f4e6c2",
   423 => x"31c849bf",
   424 => x"97f3e6c2",
   425 => x"49a14abf",
   426 => x"59f2eec2",
   427 => x"bfeeeec2",
   428 => x"c731c549",
   429 => x"29c981ff",
   430 => x"59cbf3c2",
   431 => x"97f9e6c2",
   432 => x"32c84abf",
   433 => x"97f8e6c2",
   434 => x"4aa24bbf",
   435 => x"6e9266c4",
   436 => x"c7f3c282",
   437 => x"fff2c25a",
   438 => x"c278c048",
   439 => x"7248fbf2",
   440 => x"f3c278a1",
   441 => x"f2c248cb",
   442 => x"c278bfff",
   443 => x"c248cff3",
   444 => x"78bfc3f3",
   445 => x"bfeaeec2",
   446 => x"87c9c002",
   447 => x"30c44874",
   448 => x"c9c07e70",
   449 => x"c7f3c287",
   450 => x"30c448bf",
   451 => x"eec27e70",
   452 => x"786e48ee",
   453 => x"8ef848c1",
   454 => x"4c264d26",
   455 => x"4f264b26",
   456 => x"5c5b5e0e",
   457 => x"4a710e5d",
   458 => x"bfeaeec2",
   459 => x"7287cb02",
   460 => x"722bc74b",
   461 => x"9cffc14c",
   462 => x"4b7287c9",
   463 => x"4c722bc8",
   464 => x"c29cffc3",
   465 => x"83bff7f2",
   466 => x"bfd9f5c0",
   467 => x"87d902ab",
   468 => x"5bddf5c0",
   469 => x"1ee2e6c2",
   470 => x"fdf04973",
   471 => x"7086c487",
   472 => x"87c50598",
   473 => x"e6c048c0",
   474 => x"eaeec287",
   475 => x"87d202bf",
   476 => x"91c44974",
   477 => x"81e2e6c2",
   478 => x"ffcf4d69",
   479 => x"9dffffff",
   480 => x"497487cb",
   481 => x"e6c291c2",
   482 => x"699f81e2",
   483 => x"fe48754d",
   484 => x"5e0e87c6",
   485 => x"0e5d5c5b",
   486 => x"4c7186f8",
   487 => x"87c5059c",
   488 => x"c1c348c0",
   489 => x"7ea4c887",
   490 => x"78c0486e",
   491 => x"c70266d8",
   492 => x"9766d887",
   493 => x"87c505bf",
   494 => x"e9c248c0",
   495 => x"c11ec087",
   496 => x"87f9ce49",
   497 => x"4d7086c4",
   498 => x"c2c1029d",
   499 => x"f2eec287",
   500 => x"4966d84a",
   501 => x"7087f8e1",
   502 => x"f2c00298",
   503 => x"d84a7587",
   504 => x"4bcb4966",
   505 => x"7087dde2",
   506 => x"e2c00298",
   507 => x"751ec087",
   508 => x"87c7029d",
   509 => x"c048a6c8",
   510 => x"c887c578",
   511 => x"78c148a6",
   512 => x"cd4966c8",
   513 => x"86c487f7",
   514 => x"059d4d70",
   515 => x"7587fefe",
   516 => x"cfc1029d",
   517 => x"49a5dc87",
   518 => x"7869486e",
   519 => x"c449a5da",
   520 => x"a4c448a6",
   521 => x"48699f78",
   522 => x"780866c4",
   523 => x"bfeaeec2",
   524 => x"d487d202",
   525 => x"699f49a5",
   526 => x"ffffc049",
   527 => x"d0487199",
   528 => x"c27e7030",
   529 => x"6e7ec087",
   530 => x"66c44849",
   531 => x"66c480bf",
   532 => x"7cc07808",
   533 => x"c449a4cc",
   534 => x"d079bf66",
   535 => x"79c049a4",
   536 => x"87c248c1",
   537 => x"8ef848c0",
   538 => x"0e87edfa",
   539 => x"5d5c5b5e",
   540 => x"9c4c710e",
   541 => x"87cac102",
   542 => x"6949a4c8",
   543 => x"87c2c102",
   544 => x"6c4a66d0",
   545 => x"a6d48249",
   546 => x"4d66d05a",
   547 => x"e6eec2b9",
   548 => x"baff4abf",
   549 => x"99719972",
   550 => x"87e4c002",
   551 => x"6b4ba4c4",
   552 => x"87fcf949",
   553 => x"eec27b70",
   554 => x"6c49bfe2",
   555 => x"757c7181",
   556 => x"e6eec2b9",
   557 => x"baff4abf",
   558 => x"99719972",
   559 => x"87dcff05",
   560 => x"d3f97c75",
   561 => x"1e731e87",
   562 => x"029b4b71",
   563 => x"a3c887c7",
   564 => x"c5056949",
   565 => x"c048c087",
   566 => x"f2c287f7",
   567 => x"c44abffb",
   568 => x"496949a3",
   569 => x"eec289c2",
   570 => x"7191bfe2",
   571 => x"eec24aa2",
   572 => x"6b49bfe6",
   573 => x"4aa27199",
   574 => x"5addf5c0",
   575 => x"721e66c8",
   576 => x"87d6ea49",
   577 => x"987086c4",
   578 => x"c087c405",
   579 => x"c187c248",
   580 => x"87c8f848",
   581 => x"5c5b5e0e",
   582 => x"711e0e5d",
   583 => x"4c66d44b",
   584 => x"9b732cc9",
   585 => x"87cfc102",
   586 => x"6949a3c8",
   587 => x"87c7c102",
   588 => x"d44da3d0",
   589 => x"eec27d66",
   590 => x"ff49bfe6",
   591 => x"994a6bb9",
   592 => x"03ac717e",
   593 => x"7bc087cd",
   594 => x"4aa3cc7d",
   595 => x"6a49a3c4",
   596 => x"7287c279",
   597 => x"029c748c",
   598 => x"1e4987dd",
   599 => x"cafc4973",
   600 => x"d486c487",
   601 => x"ffc74966",
   602 => x"87cb0299",
   603 => x"1ee2e6c2",
   604 => x"d0fd4973",
   605 => x"2686c487",
   606 => x"0e87ddf6",
   607 => x"5d5c5b5e",
   608 => x"d086f00e",
   609 => x"e4c059a6",
   610 => x"66cc4b66",
   611 => x"4887ca02",
   612 => x"7e7080c8",
   613 => x"c505bf6e",
   614 => x"c348c087",
   615 => x"66cc87ec",
   616 => x"7384d04c",
   617 => x"48a6c449",
   618 => x"66c4786c",
   619 => x"6e80c481",
   620 => x"66c878bf",
   621 => x"87c606a9",
   622 => x"8966c449",
   623 => x"b7c04b71",
   624 => x"87c401ab",
   625 => x"87c2c348",
   626 => x"c74866c4",
   627 => x"7e7098ff",
   628 => x"c9c1026e",
   629 => x"49c0c887",
   630 => x"4a71896e",
   631 => x"4de2e6c2",
   632 => x"b773856e",
   633 => x"87c106aa",
   634 => x"4849724a",
   635 => x"708066c4",
   636 => x"498b727c",
   637 => x"99718ac1",
   638 => x"c087d902",
   639 => x"154866e0",
   640 => x"66e0c050",
   641 => x"c080c148",
   642 => x"7258a6e4",
   643 => x"718ac149",
   644 => x"87e70599",
   645 => x"66d01ec1",
   646 => x"87cff949",
   647 => x"b7c086c4",
   648 => x"e3c106ab",
   649 => x"66e0c087",
   650 => x"b7ffc74d",
   651 => x"e2c006ab",
   652 => x"d01e7587",
   653 => x"ccfa4966",
   654 => x"85c0c887",
   655 => x"c0c8486c",
   656 => x"c87c7080",
   657 => x"1ec18bc0",
   658 => x"f84966d4",
   659 => x"86c887dd",
   660 => x"c287eec0",
   661 => x"d01ee2e6",
   662 => x"e8f94966",
   663 => x"c286c487",
   664 => x"734ae2e6",
   665 => x"806c4849",
   666 => x"49737c70",
   667 => x"99718bc1",
   668 => x"1287ce02",
   669 => x"85c17d97",
   670 => x"8bc14973",
   671 => x"f2059971",
   672 => x"abb7c087",
   673 => x"87e1fe01",
   674 => x"8ef048c1",
   675 => x"0e87c9f2",
   676 => x"5d5c5b5e",
   677 => x"9b4b710e",
   678 => x"c887c702",
   679 => x"056d4da3",
   680 => x"48ff87c5",
   681 => x"d087fdc0",
   682 => x"496c4ca3",
   683 => x"0599ffc7",
   684 => x"026c87d8",
   685 => x"1ec187c9",
   686 => x"eef64973",
   687 => x"c286c487",
   688 => x"731ee2e6",
   689 => x"87fdf749",
   690 => x"4a6c86c4",
   691 => x"c404aa6d",
   692 => x"cf48ff87",
   693 => x"7ca2c187",
   694 => x"ffc74972",
   695 => x"e2e6c299",
   696 => x"48699781",
   697 => x"1e87f1f0",
   698 => x"4b711e73",
   699 => x"e4c0029b",
   700 => x"cff3c287",
   701 => x"c24a735b",
   702 => x"e2eec28a",
   703 => x"c29249bf",
   704 => x"48bffbf2",
   705 => x"f3c28072",
   706 => x"487158d3",
   707 => x"eec230c4",
   708 => x"edc058f2",
   709 => x"cbf3c287",
   710 => x"fff2c248",
   711 => x"f3c278bf",
   712 => x"f3c248cf",
   713 => x"c278bfc3",
   714 => x"02bfeaee",
   715 => x"eec287c9",
   716 => x"c449bfe2",
   717 => x"c287c731",
   718 => x"49bfc7f3",
   719 => x"eec231c4",
   720 => x"d7ef59f2",
   721 => x"5b5e0e87",
   722 => x"4a710e5c",
   723 => x"9a724bc0",
   724 => x"87e1c002",
   725 => x"9f49a2da",
   726 => x"eec24b69",
   727 => x"cf02bfea",
   728 => x"49a2d487",
   729 => x"4c49699f",
   730 => x"9cffffc0",
   731 => x"87c234d0",
   732 => x"49744cc0",
   733 => x"fd4973b3",
   734 => x"ddee87ed",
   735 => x"5b5e0e87",
   736 => x"f40e5d5c",
   737 => x"c04a7186",
   738 => x"029a727e",
   739 => x"e6c287d8",
   740 => x"78c048de",
   741 => x"48d6e6c2",
   742 => x"bfcff3c2",
   743 => x"dae6c278",
   744 => x"cbf3c248",
   745 => x"eec278bf",
   746 => x"50c048ff",
   747 => x"bfeeeec2",
   748 => x"dee6c249",
   749 => x"aa714abf",
   750 => x"87cac403",
   751 => x"99cf4972",
   752 => x"87eac005",
   753 => x"48d9f5c0",
   754 => x"bfd6e6c2",
   755 => x"e2e6c278",
   756 => x"d6e6c21e",
   757 => x"e6c249bf",
   758 => x"a1c148d6",
   759 => x"deff7178",
   760 => x"86c487f8",
   761 => x"48d5f5c0",
   762 => x"78e2e6c2",
   763 => x"f5c087cc",
   764 => x"c048bfd5",
   765 => x"f5c080e0",
   766 => x"e6c258d9",
   767 => x"c148bfde",
   768 => x"e2e6c280",
   769 => x"0d552758",
   770 => x"97bf0000",
   771 => x"029d4dbf",
   772 => x"c387e3c2",
   773 => x"c202ade5",
   774 => x"f5c087dc",
   775 => x"cb4bbfd5",
   776 => x"4c1149a3",
   777 => x"c105accf",
   778 => x"497587d2",
   779 => x"89c199df",
   780 => x"eec291cd",
   781 => x"a3c181f2",
   782 => x"c351124a",
   783 => x"51124aa3",
   784 => x"124aa3c5",
   785 => x"4aa3c751",
   786 => x"a3c95112",
   787 => x"ce51124a",
   788 => x"51124aa3",
   789 => x"124aa3d0",
   790 => x"4aa3d251",
   791 => x"a3d45112",
   792 => x"d651124a",
   793 => x"51124aa3",
   794 => x"124aa3d8",
   795 => x"4aa3dc51",
   796 => x"a3de5112",
   797 => x"c151124a",
   798 => x"87fac07e",
   799 => x"99c84974",
   800 => x"87ebc005",
   801 => x"99d04974",
   802 => x"dc87d105",
   803 => x"cbc00266",
   804 => x"dc497387",
   805 => x"98700f66",
   806 => x"87d3c002",
   807 => x"c6c0056e",
   808 => x"f2eec287",
   809 => x"c050c048",
   810 => x"48bfd5f5",
   811 => x"c287e1c2",
   812 => x"c048ffee",
   813 => x"eec27e50",
   814 => x"c249bfee",
   815 => x"4abfdee6",
   816 => x"fb04aa71",
   817 => x"f3c287f6",
   818 => x"c005bfcf",
   819 => x"eec287c8",
   820 => x"c102bfea",
   821 => x"e6c287f8",
   822 => x"e949bfda",
   823 => x"497087c2",
   824 => x"59dee6c2",
   825 => x"c248a6c4",
   826 => x"78bfdae6",
   827 => x"bfeaeec2",
   828 => x"87d8c002",
   829 => x"cf4966c4",
   830 => x"f8ffffff",
   831 => x"c002a999",
   832 => x"4cc087c5",
   833 => x"c187e1c0",
   834 => x"87dcc04c",
   835 => x"cf4966c4",
   836 => x"a999f8ff",
   837 => x"87c8c002",
   838 => x"c048a6c8",
   839 => x"87c5c078",
   840 => x"c148a6c8",
   841 => x"4c66c878",
   842 => x"c0059c74",
   843 => x"66c487e0",
   844 => x"c289c249",
   845 => x"4abfe2ee",
   846 => x"fbf2c291",
   847 => x"e6c24abf",
   848 => x"a17248d6",
   849 => x"dee6c278",
   850 => x"f978c048",
   851 => x"48c087de",
   852 => x"c3e78ef4",
   853 => x"00000087",
   854 => x"ffffff00",
   855 => x"000d65ff",
   856 => x"000d6e00",
   857 => x"54414600",
   858 => x"20203233",
   859 => x"41460020",
   860 => x"20363154",
   861 => x"1e002020",
   862 => x"bfd4f3c2",
   863 => x"05a8dd48",
   864 => x"c3c187c9",
   865 => x"497087c8",
   866 => x"ff87c84a",
   867 => x"ffc348d4",
   868 => x"724a6878",
   869 => x"1e4f2648",
   870 => x"bfd4f3c2",
   871 => x"05a8dd48",
   872 => x"c2c187c6",
   873 => x"87d987d4",
   874 => x"c348d4ff",
   875 => x"d0ff78ff",
   876 => x"78e1c048",
   877 => x"d448d4ff",
   878 => x"d3f3c278",
   879 => x"bfd4ff48",
   880 => x"1e4f2650",
   881 => x"c048d0ff",
   882 => x"4f2678e0",
   883 => x"87e7fe1e",
   884 => x"02994970",
   885 => x"fbc087c6",
   886 => x"87f105a9",
   887 => x"4f264871",
   888 => x"5c5b5e0e",
   889 => x"c04b710e",
   890 => x"87cbfe4c",
   891 => x"02994970",
   892 => x"c087f9c0",
   893 => x"c002a9ec",
   894 => x"fbc087f2",
   895 => x"ebc002a9",
   896 => x"b766cc87",
   897 => x"87c703ac",
   898 => x"c20266d0",
   899 => x"71537187",
   900 => x"87c20299",
   901 => x"defd84c1",
   902 => x"99497087",
   903 => x"c087cd02",
   904 => x"c702a9ec",
   905 => x"a9fbc087",
   906 => x"87d5ff05",
   907 => x"c30266d0",
   908 => x"7b97c087",
   909 => x"05a9ecc0",
   910 => x"4a7487c4",
   911 => x"4a7487c5",
   912 => x"728a0ac0",
   913 => x"2687c248",
   914 => x"264c264d",
   915 => x"1e4f264b",
   916 => x"7087e4fc",
   917 => x"b7f0c049",
   918 => x"87ca04a9",
   919 => x"a9b7f9c0",
   920 => x"c087c301",
   921 => x"c1c189f0",
   922 => x"ca04a9b7",
   923 => x"b7dac187",
   924 => x"87c301a9",
   925 => x"7189f7c0",
   926 => x"0e4f2648",
   927 => x"0e5c5b5e",
   928 => x"d4ff4a71",
   929 => x"c049724c",
   930 => x"4b7087e9",
   931 => x"87c2029b",
   932 => x"d0ff8bc1",
   933 => x"c178c548",
   934 => x"49737cd5",
   935 => x"e7c131c6",
   936 => x"4abf97d0",
   937 => x"70b07148",
   938 => x"48d0ff7c",
   939 => x"487378c4",
   940 => x"0e87d6fe",
   941 => x"5d5c5b5e",
   942 => x"7186f40e",
   943 => x"48a6c44c",
   944 => x"a4c878c0",
   945 => x"bf976e7e",
   946 => x"a9c1c149",
   947 => x"c987dd05",
   948 => x"699749a4",
   949 => x"a9d2c149",
   950 => x"ca87d105",
   951 => x"699749a4",
   952 => x"a9c3c149",
   953 => x"df87c505",
   954 => x"87e1c248",
   955 => x"c087e8fa",
   956 => x"d2fec04b",
   957 => x"c049bf97",
   958 => x"87cf04a9",
   959 => x"c187cdfb",
   960 => x"d2fec083",
   961 => x"ab49bf97",
   962 => x"c087f106",
   963 => x"bf97d2fe",
   964 => x"f987cf02",
   965 => x"497087e1",
   966 => x"87c60299",
   967 => x"05a9ecc0",
   968 => x"4bc087f1",
   969 => x"7087d0f9",
   970 => x"87cbf94d",
   971 => x"f958a6cc",
   972 => x"4a7087c5",
   973 => x"976e83c1",
   974 => x"02ad49bf",
   975 => x"ffc087c7",
   976 => x"eac005ad",
   977 => x"49a4c987",
   978 => x"c8496997",
   979 => x"c702a966",
   980 => x"ffc04887",
   981 => x"87d705a8",
   982 => x"9749a4ca",
   983 => x"02aa4969",
   984 => x"ffc087c6",
   985 => x"87c705aa",
   986 => x"c148a6c4",
   987 => x"c087d378",
   988 => x"c602adec",
   989 => x"adfbc087",
   990 => x"c087c705",
   991 => x"48a6c44b",
   992 => x"66c478c1",
   993 => x"87dcfe02",
   994 => x"7387f8f8",
   995 => x"fa8ef448",
   996 => x"0e0087f5",
   997 => x"5d5c5b5e",
   998 => x"7186f80e",
   999 => x"4bd4ff4d",
  1000 => x"f3c21e75",
  1001 => x"dfff49d8",
  1002 => x"86c487e8",
  1003 => x"c4029870",
  1004 => x"e7c187fb",
  1005 => x"757ebfd2",
  1006 => x"87fffa49",
  1007 => x"c005a8de",
  1008 => x"497587eb",
  1009 => x"87e4f7c0",
  1010 => x"db029870",
  1011 => x"fcf7c287",
  1012 => x"e1c01ebf",
  1013 => x"cbf4c049",
  1014 => x"c186c487",
  1015 => x"c048d0e7",
  1016 => x"c8f8c250",
  1017 => x"87ebfe49",
  1018 => x"c2c448c1",
  1019 => x"48d0ff87",
  1020 => x"d6c178c5",
  1021 => x"754ac07b",
  1022 => x"7b1149a2",
  1023 => x"b7cb82c1",
  1024 => x"87f304aa",
  1025 => x"ffc34acc",
  1026 => x"c082c17b",
  1027 => x"04aab7e0",
  1028 => x"d0ff87f4",
  1029 => x"c378c448",
  1030 => x"78c57bff",
  1031 => x"c17bd3c1",
  1032 => x"6e78c47b",
  1033 => x"a8b7c048",
  1034 => x"87f0c206",
  1035 => x"bfe0f3c2",
  1036 => x"74486e4c",
  1037 => x"747e7088",
  1038 => x"fdc1029c",
  1039 => x"e2e6c287",
  1040 => x"48a6c44d",
  1041 => x"8c78c0c8",
  1042 => x"03acb7c0",
  1043 => x"c0c887c6",
  1044 => x"4cc078a4",
  1045 => x"97d3f3c2",
  1046 => x"99d049bf",
  1047 => x"c087d102",
  1048 => x"d8f3c21e",
  1049 => x"87dde149",
  1050 => x"497086c4",
  1051 => x"87eec04a",
  1052 => x"1ee2e6c2",
  1053 => x"49d8f3c2",
  1054 => x"c487cae1",
  1055 => x"4a497086",
  1056 => x"c848d0ff",
  1057 => x"d4c178c5",
  1058 => x"c47b157b",
  1059 => x"88c14866",
  1060 => x"7058a6c8",
  1061 => x"f0ff0598",
  1062 => x"48d0ff87",
  1063 => x"9a7278c4",
  1064 => x"c087c505",
  1065 => x"87c7c148",
  1066 => x"f3c21ec1",
  1067 => x"deff49d8",
  1068 => x"86c487f9",
  1069 => x"fe059c74",
  1070 => x"486e87c3",
  1071 => x"06a8b7c0",
  1072 => x"f3c287d1",
  1073 => x"78c048d8",
  1074 => x"78c080d0",
  1075 => x"f3c280f4",
  1076 => x"6e78bfe4",
  1077 => x"a8b7c048",
  1078 => x"87d0fd01",
  1079 => x"c548d0ff",
  1080 => x"7bd3c178",
  1081 => x"78c47bc0",
  1082 => x"c2c048c1",
  1083 => x"f848c087",
  1084 => x"264d268e",
  1085 => x"264b264c",
  1086 => x"5b5e0e4f",
  1087 => x"1e0e5d5c",
  1088 => x"4cc04b71",
  1089 => x"c004ab4d",
  1090 => x"fac087e8",
  1091 => x"9d751ef3",
  1092 => x"c087c402",
  1093 => x"c187c24a",
  1094 => x"e949724a",
  1095 => x"86c487df",
  1096 => x"84c17e70",
  1097 => x"87c2056e",
  1098 => x"85c14c73",
  1099 => x"ff06ac73",
  1100 => x"486e87d8",
  1101 => x"87f9fe26",
  1102 => x"c44a711e",
  1103 => x"87c50566",
  1104 => x"cef94972",
  1105 => x"0e4f2687",
  1106 => x"5d5c5b5e",
  1107 => x"4c711e0e",
  1108 => x"c291de49",
  1109 => x"714dc0f4",
  1110 => x"026d9785",
  1111 => x"c287dcc1",
  1112 => x"4abfecf3",
  1113 => x"49728274",
  1114 => x"7087cefe",
  1115 => x"c0026e7e",
  1116 => x"f3c287f2",
  1117 => x"4a6e4bf4",
  1118 => x"fcfe49cb",
  1119 => x"4b7487ea",
  1120 => x"e7c193cb",
  1121 => x"83c483e4",
  1122 => x"7bffc6c1",
  1123 => x"ccc14974",
  1124 => x"7b7587c7",
  1125 => x"97d1e7c1",
  1126 => x"c21e49bf",
  1127 => x"fe49f4f3",
  1128 => x"86c487d6",
  1129 => x"cbc14974",
  1130 => x"49c087ef",
  1131 => x"87cecdc1",
  1132 => x"48d4f3c2",
  1133 => x"49c178c0",
  1134 => x"2687d4dd",
  1135 => x"4c87f2fc",
  1136 => x"6964616f",
  1137 => x"2e2e676e",
  1138 => x"5e0e002e",
  1139 => x"710e5c5b",
  1140 => x"f3c24a4b",
  1141 => x"7282bfec",
  1142 => x"87ddfc49",
  1143 => x"029c4c70",
  1144 => x"e54987c4",
  1145 => x"f3c287df",
  1146 => x"78c048ec",
  1147 => x"dedc49c1",
  1148 => x"87fffb87",
  1149 => x"5c5b5e0e",
  1150 => x"86f40e5d",
  1151 => x"4de2e6c2",
  1152 => x"a6c44cc0",
  1153 => x"c278c048",
  1154 => x"49bfecf3",
  1155 => x"c106a9c0",
  1156 => x"e6c287c1",
  1157 => x"029848e2",
  1158 => x"c087f8c0",
  1159 => x"c81ef3fa",
  1160 => x"87c70266",
  1161 => x"c048a6c4",
  1162 => x"c487c578",
  1163 => x"78c148a6",
  1164 => x"e54966c4",
  1165 => x"86c487c7",
  1166 => x"84c14d70",
  1167 => x"c14866c4",
  1168 => x"58a6c880",
  1169 => x"bfecf3c2",
  1170 => x"c603ac49",
  1171 => x"059d7587",
  1172 => x"c087c8ff",
  1173 => x"029d754c",
  1174 => x"c087e0c3",
  1175 => x"c81ef3fa",
  1176 => x"87c70266",
  1177 => x"c048a6cc",
  1178 => x"cc87c578",
  1179 => x"78c148a6",
  1180 => x"e44966cc",
  1181 => x"86c487c7",
  1182 => x"026e7e70",
  1183 => x"6e87e9c2",
  1184 => x"9781cb49",
  1185 => x"99d04969",
  1186 => x"87d6c102",
  1187 => x"4acac7c1",
  1188 => x"91cb4974",
  1189 => x"81e4e7c1",
  1190 => x"81c87972",
  1191 => x"7451ffc3",
  1192 => x"c291de49",
  1193 => x"714dc0f4",
  1194 => x"97c1c285",
  1195 => x"49a5c17d",
  1196 => x"c251e0c0",
  1197 => x"bf97f2ee",
  1198 => x"c187d202",
  1199 => x"4ba5c284",
  1200 => x"4af2eec2",
  1201 => x"f7fe49db",
  1202 => x"dbc187de",
  1203 => x"49a5cd87",
  1204 => x"84c151c0",
  1205 => x"6e4ba5c2",
  1206 => x"fe49cb4a",
  1207 => x"c187c9f7",
  1208 => x"c5c187c6",
  1209 => x"49744ac7",
  1210 => x"e7c191cb",
  1211 => x"797281e4",
  1212 => x"97f2eec2",
  1213 => x"87d802bf",
  1214 => x"91de4974",
  1215 => x"f4c284c1",
  1216 => x"83714bc0",
  1217 => x"4af2eec2",
  1218 => x"f6fe49dd",
  1219 => x"87d887da",
  1220 => x"93de4b74",
  1221 => x"83c0f4c2",
  1222 => x"c049a3cb",
  1223 => x"7384c151",
  1224 => x"49cb4a6e",
  1225 => x"87c0f6fe",
  1226 => x"c14866c4",
  1227 => x"58a6c880",
  1228 => x"c003acc7",
  1229 => x"056e87c5",
  1230 => x"7487e0fc",
  1231 => x"f68ef448",
  1232 => x"731e87ef",
  1233 => x"494b711e",
  1234 => x"e7c191cb",
  1235 => x"a1c881e4",
  1236 => x"d0e7c14a",
  1237 => x"c9501248",
  1238 => x"fec04aa1",
  1239 => x"501248d2",
  1240 => x"e7c181ca",
  1241 => x"501148d1",
  1242 => x"97d1e7c1",
  1243 => x"c01e49bf",
  1244 => x"87c4f749",
  1245 => x"48d4f3c2",
  1246 => x"49c178de",
  1247 => x"2687d0d6",
  1248 => x"1e87f2f5",
  1249 => x"cb494a71",
  1250 => x"e4e7c191",
  1251 => x"1181c881",
  1252 => x"d8f3c248",
  1253 => x"ecf3c258",
  1254 => x"c178c048",
  1255 => x"87efd549",
  1256 => x"c01e4f26",
  1257 => x"d5c5c149",
  1258 => x"1e4f2687",
  1259 => x"d2029971",
  1260 => x"f9e8c187",
  1261 => x"f750c048",
  1262 => x"c3cec180",
  1263 => x"dde7c140",
  1264 => x"c187ce78",
  1265 => x"c148f5e8",
  1266 => x"fc78d6e7",
  1267 => x"e2cec180",
  1268 => x"0e4f2678",
  1269 => x"0e5c5b5e",
  1270 => x"cb4a4c71",
  1271 => x"e4e7c192",
  1272 => x"49a2c882",
  1273 => x"974ba2c9",
  1274 => x"971e4b6b",
  1275 => x"ca1e4969",
  1276 => x"c0491282",
  1277 => x"c087f5e5",
  1278 => x"87d3d449",
  1279 => x"c2c14974",
  1280 => x"8ef887d7",
  1281 => x"1e87ecf3",
  1282 => x"4b711e73",
  1283 => x"87c3ff49",
  1284 => x"fefe4973",
  1285 => x"87ddf387",
  1286 => x"711e731e",
  1287 => x"4aa3c64b",
  1288 => x"c187db02",
  1289 => x"87d6028a",
  1290 => x"dac1028a",
  1291 => x"c0028a87",
  1292 => x"028a87fc",
  1293 => x"8a87e1c0",
  1294 => x"c187cb02",
  1295 => x"49c787db",
  1296 => x"c187c0fd",
  1297 => x"f3c287de",
  1298 => x"c102bfec",
  1299 => x"c14887cb",
  1300 => x"f0f3c288",
  1301 => x"87c1c158",
  1302 => x"bff0f3c2",
  1303 => x"87f9c002",
  1304 => x"bfecf3c2",
  1305 => x"c280c148",
  1306 => x"c058f0f3",
  1307 => x"f3c287eb",
  1308 => x"c649bfec",
  1309 => x"f0f3c289",
  1310 => x"a9b7c059",
  1311 => x"c287da03",
  1312 => x"c048ecf3",
  1313 => x"c287d278",
  1314 => x"02bff0f3",
  1315 => x"f3c287cb",
  1316 => x"c648bfec",
  1317 => x"f0f3c280",
  1318 => x"d149c058",
  1319 => x"497387f1",
  1320 => x"87f5ffc0",
  1321 => x"1e87cef1",
  1322 => x"4b711e73",
  1323 => x"48d4f3c2",
  1324 => x"49c078dd",
  1325 => x"7387d8d1",
  1326 => x"dcffc049",
  1327 => x"87f5f087",
  1328 => x"5c5b5e0e",
  1329 => x"cc4c710e",
  1330 => x"4b741e66",
  1331 => x"e7c193cb",
  1332 => x"a3c483e4",
  1333 => x"fe496a4a",
  1334 => x"c187ddef",
  1335 => x"c87bc2cd",
  1336 => x"66d449a3",
  1337 => x"49a3c951",
  1338 => x"ca5166d8",
  1339 => x"66dc49a3",
  1340 => x"feef2651",
  1341 => x"5b5e0e87",
  1342 => x"ff0e5d5c",
  1343 => x"a6dc86cc",
  1344 => x"48a6c859",
  1345 => x"80c478c0",
  1346 => x"7866c8c1",
  1347 => x"78c180c4",
  1348 => x"78c180c4",
  1349 => x"48f0f3c2",
  1350 => x"f3c278c1",
  1351 => x"de48bfd4",
  1352 => x"87cb05a8",
  1353 => x"7087cdf3",
  1354 => x"59a6cc49",
  1355 => x"e187dbce",
  1356 => x"d7e287e5",
  1357 => x"87ffe087",
  1358 => x"fbc04c70",
  1359 => x"ddc102ac",
  1360 => x"0566d887",
  1361 => x"c087cfc1",
  1362 => x"1ec11e1e",
  1363 => x"1ec7e9c1",
  1364 => x"ebfd49c0",
  1365 => x"c186d087",
  1366 => x"c44866c4",
  1367 => x"6e7e7080",
  1368 => x"81c749bf",
  1369 => x"fbc05174",
  1370 => x"87cf02ac",
  1371 => x"1ed81ec1",
  1372 => x"49bf66c8",
  1373 => x"e7e181c8",
  1374 => x"c186c887",
  1375 => x"c04866c8",
  1376 => x"87c701a8",
  1377 => x"c148a6c8",
  1378 => x"c187ce78",
  1379 => x"c14866c8",
  1380 => x"58a6d088",
  1381 => x"f3e087c3",
  1382 => x"48a6d087",
  1383 => x"9c7478c2",
  1384 => x"87e2cc02",
  1385 => x"c14866c8",
  1386 => x"03a866cc",
  1387 => x"c487d7cc",
  1388 => x"78c048a6",
  1389 => x"78c080d8",
  1390 => x"87fbdeff",
  1391 => x"66d84c70",
  1392 => x"05a8dd48",
  1393 => x"a6dc87c6",
  1394 => x"7866d848",
  1395 => x"05acd0c1",
  1396 => x"ff87ebc0",
  1397 => x"ff87e0de",
  1398 => x"7087dcde",
  1399 => x"acecc04c",
  1400 => x"ff87c605",
  1401 => x"7087e5df",
  1402 => x"acd0c14c",
  1403 => x"d487c805",
  1404 => x"80c14866",
  1405 => x"c158a6d8",
  1406 => x"ff02acd0",
  1407 => x"e0c087d5",
  1408 => x"66d848a6",
  1409 => x"4866dc78",
  1410 => x"a866e0c0",
  1411 => x"87c8ca05",
  1412 => x"48a6e4c0",
  1413 => x"80c478c0",
  1414 => x"4d7478c0",
  1415 => x"028dfbc0",
  1416 => x"c987cec9",
  1417 => x"87db028d",
  1418 => x"c1028dc2",
  1419 => x"8dc987f7",
  1420 => x"87d1c402",
  1421 => x"c1028dc4",
  1422 => x"8dc187c2",
  1423 => x"87c5c402",
  1424 => x"c887e8c8",
  1425 => x"91cb4966",
  1426 => x"8166c4c1",
  1427 => x"6a4aa1c4",
  1428 => x"c11e717e",
  1429 => x"c448c2e4",
  1430 => x"a1cc4966",
  1431 => x"7141204a",
  1432 => x"f8ff05aa",
  1433 => x"26511087",
  1434 => x"e7d2c149",
  1435 => x"dbddff79",
  1436 => x"c04c7087",
  1437 => x"c148a6e8",
  1438 => x"87f5c778",
  1439 => x"c048a6c4",
  1440 => x"dbff78f0",
  1441 => x"4c7087f1",
  1442 => x"02acecc0",
  1443 => x"c887c3c0",
  1444 => x"ecc05ca6",
  1445 => x"87cd02ac",
  1446 => x"87dbdbff",
  1447 => x"ecc04c70",
  1448 => x"f3ff05ac",
  1449 => x"acecc087",
  1450 => x"87c4c002",
  1451 => x"87c7dbff",
  1452 => x"d81e66c4",
  1453 => x"d81e4966",
  1454 => x"c11e4966",
  1455 => x"d81ec7e9",
  1456 => x"fbf74966",
  1457 => x"ca1ec087",
  1458 => x"66e0c01e",
  1459 => x"c191cb49",
  1460 => x"d88166dc",
  1461 => x"a1c448a6",
  1462 => x"bf66d878",
  1463 => x"ffdbff49",
  1464 => x"c086d887",
  1465 => x"c106a8b7",
  1466 => x"1ec187cb",
  1467 => x"66c81ede",
  1468 => x"dbff49bf",
  1469 => x"86c887ea",
  1470 => x"c0484970",
  1471 => x"ecc08808",
  1472 => x"b7c058a6",
  1473 => x"ecc006a8",
  1474 => x"66e8c087",
  1475 => x"a8b7dd48",
  1476 => x"87e1c003",
  1477 => x"c049bf6e",
  1478 => x"c08166e8",
  1479 => x"e8c051e0",
  1480 => x"81c14966",
  1481 => x"c281bf6e",
  1482 => x"e8c051c1",
  1483 => x"81c24966",
  1484 => x"c081bf6e",
  1485 => x"4866d051",
  1486 => x"a6d480c1",
  1487 => x"80d84858",
  1488 => x"ecc478c1",
  1489 => x"c6dcff87",
  1490 => x"a6ecc087",
  1491 => x"fedbff58",
  1492 => x"a6f0c087",
  1493 => x"a8ecc058",
  1494 => x"87c9c005",
  1495 => x"e8c048a6",
  1496 => x"c4c07866",
  1497 => x"ced8ff87",
  1498 => x"4966c887",
  1499 => x"c4c191cb",
  1500 => x"80714866",
  1501 => x"c458a6c8",
  1502 => x"82c84a66",
  1503 => x"ca4966c4",
  1504 => x"66e8c081",
  1505 => x"66ecc051",
  1506 => x"c081c149",
  1507 => x"c18966e8",
  1508 => x"70307148",
  1509 => x"7189c149",
  1510 => x"f7c27a97",
  1511 => x"c049bfdc",
  1512 => x"972966e8",
  1513 => x"71484a6a",
  1514 => x"a6f4c098",
  1515 => x"4966c458",
  1516 => x"7e6981c4",
  1517 => x"4866e0c0",
  1518 => x"02a866dc",
  1519 => x"dc87c8c0",
  1520 => x"78c048a6",
  1521 => x"dc87c5c0",
  1522 => x"78c148a6",
  1523 => x"c01e66dc",
  1524 => x"66c81ee0",
  1525 => x"c7d8ff49",
  1526 => x"7086c887",
  1527 => x"acb7c04c",
  1528 => x"87d6c106",
  1529 => x"8074486e",
  1530 => x"e0c07e70",
  1531 => x"6e897449",
  1532 => x"ffe3c14b",
  1533 => x"e2fe714a",
  1534 => x"486e87ee",
  1535 => x"7e7080c2",
  1536 => x"4866e4c0",
  1537 => x"e8c080c1",
  1538 => x"f0c058a6",
  1539 => x"81c14966",
  1540 => x"c002a970",
  1541 => x"4dc087c5",
  1542 => x"c187c2c0",
  1543 => x"c21e754d",
  1544 => x"e0c049a4",
  1545 => x"70887148",
  1546 => x"66c81e49",
  1547 => x"efd6ff49",
  1548 => x"c086c887",
  1549 => x"ff01a8b7",
  1550 => x"e4c087c6",
  1551 => x"d3c00266",
  1552 => x"4966c487",
  1553 => x"e4c081c9",
  1554 => x"66c45166",
  1555 => x"d3cfc148",
  1556 => x"87cec078",
  1557 => x"c94966c4",
  1558 => x"c451c281",
  1559 => x"d0c14866",
  1560 => x"e8c078c7",
  1561 => x"78c148a6",
  1562 => x"ff87c6c0",
  1563 => x"7087ddd5",
  1564 => x"66e8c04c",
  1565 => x"87f5c002",
  1566 => x"cc4866c8",
  1567 => x"c004a866",
  1568 => x"66c887cb",
  1569 => x"cc80c148",
  1570 => x"e0c058a6",
  1571 => x"4866cc87",
  1572 => x"a6d088c1",
  1573 => x"87d5c058",
  1574 => x"05acc6c1",
  1575 => x"d087c8c0",
  1576 => x"80c14866",
  1577 => x"ff58a6d4",
  1578 => x"7087e1d4",
  1579 => x"4866d44c",
  1580 => x"a6d880c1",
  1581 => x"029c7458",
  1582 => x"c887cbc0",
  1583 => x"ccc14866",
  1584 => x"f304a866",
  1585 => x"d3ff87e9",
  1586 => x"66c887f9",
  1587 => x"03a8c748",
  1588 => x"c287e5c0",
  1589 => x"c048f0f3",
  1590 => x"4966c878",
  1591 => x"c4c191cb",
  1592 => x"a1c48166",
  1593 => x"c04a6a4a",
  1594 => x"66c87952",
  1595 => x"cc80c148",
  1596 => x"a8c758a6",
  1597 => x"87dbff04",
  1598 => x"ff8eccff",
  1599 => x"3a87f2df",
  1600 => x"49440020",
  1601 => x"77532050",
  1602 => x"68637469",
  1603 => x"1e007365",
  1604 => x"4b711e73",
  1605 => x"87c6029b",
  1606 => x"48ecf3c2",
  1607 => x"1ec778c0",
  1608 => x"bfecf3c2",
  1609 => x"e7c11e49",
  1610 => x"f3c21ee4",
  1611 => x"ef49bfd4",
  1612 => x"86cc87c3",
  1613 => x"bfd4f3c2",
  1614 => x"87efe949",
  1615 => x"c8029b73",
  1616 => x"e4e7c187",
  1617 => x"e2eec049",
  1618 => x"e8deff87",
  1619 => x"d5c71e87",
  1620 => x"fe49c187",
  1621 => x"e5fe87f9",
  1622 => x"987087e9",
  1623 => x"fe87cd02",
  1624 => x"7087c2ed",
  1625 => x"87c40298",
  1626 => x"87c24ac1",
  1627 => x"9a724ac0",
  1628 => x"c087ce05",
  1629 => x"e2e6c11e",
  1630 => x"ccfac049",
  1631 => x"fe86c487",
  1632 => x"effcc087",
  1633 => x"c11ec087",
  1634 => x"c049ede6",
  1635 => x"c087faf9",
  1636 => x"f5fec01e",
  1637 => x"c0497087",
  1638 => x"c387eef9",
  1639 => x"8ef887c7",
  1640 => x"44534f26",
  1641 => x"69616620",
  1642 => x"2e64656c",
  1643 => x"6f6f4200",
  1644 => x"676e6974",
  1645 => x"002e2e2e",
  1646 => x"ecf3c21e",
  1647 => x"c278c048",
  1648 => x"c048d4f3",
  1649 => x"87c5fe78",
  1650 => x"87ddfec0",
  1651 => x"4f2648c0",
  1652 => x"00010000",
  1653 => x"20800000",
  1654 => x"74697845",
  1655 => x"42208000",
  1656 => x"006b6361",
  1657 => x"00001383",
  1658 => x"00002d00",
  1659 => x"83000000",
  1660 => x"1e000013",
  1661 => x"0000002d",
  1662 => x"13830000",
  1663 => x"2d3c0000",
  1664 => x"00000000",
  1665 => x"00138300",
  1666 => x"002d5a00",
  1667 => x"00000000",
  1668 => x"00001383",
  1669 => x"00002d78",
  1670 => x"83000000",
  1671 => x"96000013",
  1672 => x"0000002d",
  1673 => x"13830000",
  1674 => x"2db40000",
  1675 => x"00000000",
  1676 => x"00138300",
  1677 => x"00000000",
  1678 => x"00000000",
  1679 => x"00001418",
  1680 => x"00000000",
  1681 => x"4c000000",
  1682 => x"2064616f",
  1683 => x"1e002e2a",
  1684 => x"c048f0fe",
  1685 => x"7909cd78",
  1686 => x"1e4f2609",
  1687 => x"bff0fe1e",
  1688 => x"2626487e",
  1689 => x"f0fe1e4f",
  1690 => x"2678c148",
  1691 => x"f0fe1e4f",
  1692 => x"2678c048",
  1693 => x"4a711e4f",
  1694 => x"265252c0",
  1695 => x"5b5e0e4f",
  1696 => x"f40e5d5c",
  1697 => x"974d7186",
  1698 => x"a5c17e6d",
  1699 => x"486c974c",
  1700 => x"6e58a6c8",
  1701 => x"a866c448",
  1702 => x"ff87c505",
  1703 => x"87e6c048",
  1704 => x"c287caff",
  1705 => x"6c9749a5",
  1706 => x"4ba3714b",
  1707 => x"974b6b97",
  1708 => x"486e7e6c",
  1709 => x"a6c880c1",
  1710 => x"cc98c758",
  1711 => x"977058a6",
  1712 => x"87e1fe7c",
  1713 => x"8ef44873",
  1714 => x"4c264d26",
  1715 => x"4f264b26",
  1716 => x"5c5b5e0e",
  1717 => x"7186f40e",
  1718 => x"4a66d84c",
  1719 => x"c29affc3",
  1720 => x"6c974ba4",
  1721 => x"49a17349",
  1722 => x"6c975172",
  1723 => x"c1486e7e",
  1724 => x"58a6c880",
  1725 => x"a6cc98c7",
  1726 => x"f4547058",
  1727 => x"87caff8e",
  1728 => x"e8fd1e1e",
  1729 => x"4abfe087",
  1730 => x"c0e0c049",
  1731 => x"87cb0299",
  1732 => x"f7c21e72",
  1733 => x"f7fe49d2",
  1734 => x"fc86c487",
  1735 => x"7e7087fd",
  1736 => x"2687c2fd",
  1737 => x"c21e4f26",
  1738 => x"fd49d2f7",
  1739 => x"ecc187c7",
  1740 => x"dafc49c0",
  1741 => x"87c7c487",
  1742 => x"ff1e4f26",
  1743 => x"e1c848d0",
  1744 => x"48d4ff78",
  1745 => x"66c478c5",
  1746 => x"c387c302",
  1747 => x"66c878e0",
  1748 => x"ff87c602",
  1749 => x"f0c348d4",
  1750 => x"48d4ff78",
  1751 => x"d0ff7871",
  1752 => x"78e1c848",
  1753 => x"2678e0c0",
  1754 => x"5b5e0e4f",
  1755 => x"4c710e5c",
  1756 => x"49d2f7c2",
  1757 => x"7087c6fc",
  1758 => x"aab7c04a",
  1759 => x"87e2c204",
  1760 => x"05aaf0c3",
  1761 => x"f0c187c9",
  1762 => x"78c148ee",
  1763 => x"c387c3c2",
  1764 => x"c905aae0",
  1765 => x"f2f0c187",
  1766 => x"c178c148",
  1767 => x"f0c187f4",
  1768 => x"c602bff2",
  1769 => x"a2c0c287",
  1770 => x"7287c24b",
  1771 => x"059c744b",
  1772 => x"f0c187d1",
  1773 => x"c11ebfee",
  1774 => x"1ebff2f0",
  1775 => x"f9fd4972",
  1776 => x"c186c887",
  1777 => x"02bfeef0",
  1778 => x"7387e0c0",
  1779 => x"29b7c449",
  1780 => x"cef2c191",
  1781 => x"cf4a7381",
  1782 => x"c192c29a",
  1783 => x"70307248",
  1784 => x"72baff4a",
  1785 => x"70986948",
  1786 => x"7387db79",
  1787 => x"29b7c449",
  1788 => x"cef2c191",
  1789 => x"cf4a7381",
  1790 => x"c392c29a",
  1791 => x"70307248",
  1792 => x"b069484a",
  1793 => x"f0c17970",
  1794 => x"78c048f2",
  1795 => x"48eef0c1",
  1796 => x"f7c278c0",
  1797 => x"e4f949d2",
  1798 => x"c04a7087",
  1799 => x"fd03aab7",
  1800 => x"48c087de",
  1801 => x"4d2687c2",
  1802 => x"4b264c26",
  1803 => x"00004f26",
  1804 => x"00000000",
  1805 => x"711e0000",
  1806 => x"ecfc494a",
  1807 => x"1e4f2687",
  1808 => x"49724ac0",
  1809 => x"f2c191c4",
  1810 => x"79c081ce",
  1811 => x"b7d082c1",
  1812 => x"87ee04aa",
  1813 => x"5e0e4f26",
  1814 => x"0e5d5c5b",
  1815 => x"ccf84d71",
  1816 => x"c44a7587",
  1817 => x"c1922ab7",
  1818 => x"7582cef2",
  1819 => x"c29ccf4c",
  1820 => x"4b496a94",
  1821 => x"9bc32b74",
  1822 => x"307448c2",
  1823 => x"bcff4c70",
  1824 => x"98714874",
  1825 => x"dcf77a70",
  1826 => x"fe487387",
  1827 => x"000087d8",
  1828 => x"00000000",
  1829 => x"00000000",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00000000",
  1834 => x"00000000",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"00000000",
  1842 => x"00000000",
  1843 => x"ff1e0000",
  1844 => x"e1c848d0",
  1845 => x"ff487178",
  1846 => x"c47808d4",
  1847 => x"d4ff4866",
  1848 => x"4f267808",
  1849 => x"c44a711e",
  1850 => x"721e4966",
  1851 => x"87deff49",
  1852 => x"c048d0ff",
  1853 => x"262678e0",
  1854 => x"1e731e4f",
  1855 => x"66c84b71",
  1856 => x"4a731e49",
  1857 => x"49a2e0c1",
  1858 => x"2687d9ff",
  1859 => x"4d2687c4",
  1860 => x"4b264c26",
  1861 => x"731e4f26",
  1862 => x"4b4a711e",
  1863 => x"03abb7c2",
  1864 => x"49a387c8",
  1865 => x"9affc34a",
  1866 => x"a3ce87c7",
  1867 => x"ffc34a49",
  1868 => x"4966c89a",
  1869 => x"fe49721e",
  1870 => x"ff2687ea",
  1871 => x"ff1e87d4",
  1872 => x"ffc34ad4",
  1873 => x"48d0ff7a",
  1874 => x"de78e1c0",
  1875 => x"dcf7c27a",
  1876 => x"48497abf",
  1877 => x"7a7028c8",
  1878 => x"28d04871",
  1879 => x"48717a70",
  1880 => x"7a7028d8",
  1881 => x"c048d0ff",
  1882 => x"4f2678e0",
  1883 => x"5c5b5e0e",
  1884 => x"4c710e5d",
  1885 => x"bfdcf7c2",
  1886 => x"2b744b4d",
  1887 => x"c19b66d0",
  1888 => x"ab66d483",
  1889 => x"c087c204",
  1890 => x"d04a744b",
  1891 => x"31724966",
  1892 => x"9975b9ff",
  1893 => x"30724873",
  1894 => x"71484a70",
  1895 => x"e0f7c2b0",
  1896 => x"87dafe58",
  1897 => x"4c264d26",
  1898 => x"4f264b26",
  1899 => x"5c5b5e0e",
  1900 => x"711e0e5d",
  1901 => x"e0f7c24c",
  1902 => x"c04ac04b",
  1903 => x"ccfe49f4",
  1904 => x"1e7487c3",
  1905 => x"49e0f7c2",
  1906 => x"87c6e7fe",
  1907 => x"497086c4",
  1908 => x"eac00299",
  1909 => x"a61ec487",
  1910 => x"f7c21e4d",
  1911 => x"eefe49e0",
  1912 => x"86c887d9",
  1913 => x"d6029870",
  1914 => x"c14a7587",
  1915 => x"c449f5f8",
  1916 => x"f5c9fe4b",
  1917 => x"02987087",
  1918 => x"48c087ca",
  1919 => x"c087edc0",
  1920 => x"87e8c048",
  1921 => x"c187f3c0",
  1922 => x"987087c4",
  1923 => x"c087c802",
  1924 => x"987087fc",
  1925 => x"c287f805",
  1926 => x"02bfc0f8",
  1927 => x"f7c287cc",
  1928 => x"f8c248dc",
  1929 => x"fc78bfc0",
  1930 => x"48c187d4",
  1931 => x"264d2626",
  1932 => x"264b264c",
  1933 => x"52415b4f",
  1934 => x"c01e0043",
  1935 => x"e0f7c21e",
  1936 => x"cfebfe49",
  1937 => x"f8f7c287",
  1938 => x"2678c048",
  1939 => x"5e0e4f26",
  1940 => x"0e5d5c5b",
  1941 => x"a6c486f4",
  1942 => x"c278c048",
  1943 => x"48bff8f7",
  1944 => x"03a8b7c3",
  1945 => x"f7c287d1",
  1946 => x"c148bff8",
  1947 => x"fcf7c280",
  1948 => x"48fbc058",
  1949 => x"c287e2c6",
  1950 => x"fe49e0f7",
  1951 => x"7087d0f0",
  1952 => x"f8f7c24c",
  1953 => x"8ac34abf",
  1954 => x"c187d802",
  1955 => x"cbc5028a",
  1956 => x"c2028a87",
  1957 => x"028a87f6",
  1958 => x"8a87cdc1",
  1959 => x"87e2c302",
  1960 => x"c087e1c5",
  1961 => x"c44a754d",
  1962 => x"f7c0c292",
  1963 => x"f4f7c282",
  1964 => x"70807548",
  1965 => x"bf976e7e",
  1966 => x"6e4b494b",
  1967 => x"50a3c148",
  1968 => x"4811816a",
  1969 => x"7058a6cc",
  1970 => x"87c402ac",
  1971 => x"50c0486e",
  1972 => x"c70566c8",
  1973 => x"f8f7c287",
  1974 => x"78a5c448",
  1975 => x"b7c485c1",
  1976 => x"c0ff04ad",
  1977 => x"87dcc487",
  1978 => x"bfc4f8c2",
  1979 => x"a8b7c848",
  1980 => x"ca87d101",
  1981 => x"87cc02ac",
  1982 => x"c702accd",
  1983 => x"acb7c087",
  1984 => x"87f3c003",
  1985 => x"bfc4f8c2",
  1986 => x"abb7c84b",
  1987 => x"c287d203",
  1988 => x"7349c8f8",
  1989 => x"51e0c081",
  1990 => x"b7c883c1",
  1991 => x"eeff04ab",
  1992 => x"d0f8c287",
  1993 => x"50d2c148",
  1994 => x"c150cfc1",
  1995 => x"50c050cd",
  1996 => x"78c380e4",
  1997 => x"c287cdc3",
  1998 => x"49bfc4f8",
  1999 => x"c280c148",
  2000 => x"4858c8f8",
  2001 => x"7481a0c4",
  2002 => x"87f8c251",
  2003 => x"acb7f0c0",
  2004 => x"c087da04",
  2005 => x"01acb7f9",
  2006 => x"f7c287d3",
  2007 => x"ca49bffc",
  2008 => x"c04a7491",
  2009 => x"f7c28af0",
  2010 => x"a17248fc",
  2011 => x"02acca78",
  2012 => x"cd87c6c0",
  2013 => x"cbc205ac",
  2014 => x"f8f7c287",
  2015 => x"c278c348",
  2016 => x"f0c087c2",
  2017 => x"db04acb7",
  2018 => x"b7f9c087",
  2019 => x"d3c001ac",
  2020 => x"c0f8c287",
  2021 => x"91d049bf",
  2022 => x"f0c04a74",
  2023 => x"c0f8c28a",
  2024 => x"78a17248",
  2025 => x"acb7c1c1",
  2026 => x"87dbc004",
  2027 => x"acb7c6c1",
  2028 => x"87d3c001",
  2029 => x"bfc0f8c2",
  2030 => x"7491d049",
  2031 => x"8af7c04a",
  2032 => x"48c0f8c2",
  2033 => x"ca78a172",
  2034 => x"c6c002ac",
  2035 => x"05accd87",
  2036 => x"c287f1c0",
  2037 => x"c348f8f7",
  2038 => x"87e8c078",
  2039 => x"05ace2c0",
  2040 => x"c487c9c0",
  2041 => x"fbc048a6",
  2042 => x"87d8c078",
  2043 => x"c002acca",
  2044 => x"accd87c6",
  2045 => x"87c9c005",
  2046 => x"48f8f7c2",
  2047 => x"c3c078c3",
  2048 => x"5ca6c887",
  2049 => x"03acb7c0",
  2050 => x"4887c4c0",
  2051 => x"c487cac0",
  2052 => x"c6f90266",
  2053 => x"ffc34887",
  2054 => x"f88ef499",
  2055 => x"4f4387cf",
  2056 => x"003d464e",
  2057 => x"00444f4d",
  2058 => x"454d414e",
  2059 => x"46454400",
  2060 => x"544c5541",
  2061 => x"1e00303d",
  2062 => x"24000020",
  2063 => x"28000020",
  2064 => x"2d000020",
  2065 => x"1e000020",
  2066 => x"c848d0ff",
  2067 => x"487178c9",
  2068 => x"7808d4ff",
  2069 => x"711e4f26",
  2070 => x"87eb494a",
  2071 => x"c848d0ff",
  2072 => x"1e4f2678",
  2073 => x"4b711e73",
  2074 => x"bfe0f8c2",
  2075 => x"c287c302",
  2076 => x"d0ff87eb",
  2077 => x"78c9c848",
  2078 => x"e0c04973",
  2079 => x"48d4ffb1",
  2080 => x"f8c27871",
  2081 => x"78c048d4",
  2082 => x"c50266c8",
  2083 => x"49ffc387",
  2084 => x"49c087c2",
  2085 => x"59dcf8c2",
  2086 => x"c60266cc",
  2087 => x"d5d5c587",
  2088 => x"cf87c44a",
  2089 => x"c24affff",
  2090 => x"c25ae0f8",
  2091 => x"c148e0f8",
  2092 => x"2687c478",
  2093 => x"264c264d",
  2094 => x"0e4f264b",
  2095 => x"5d5c5b5e",
  2096 => x"c24a710e",
  2097 => x"4cbfdcf8",
  2098 => x"cb029a72",
  2099 => x"91c84987",
  2100 => x"4bd9c1c2",
  2101 => x"87c48371",
  2102 => x"4bd9c5c2",
  2103 => x"49134dc0",
  2104 => x"f8c29974",
  2105 => x"ffb9bfd8",
  2106 => x"787148d4",
  2107 => x"852cb7c1",
  2108 => x"04adb7c8",
  2109 => x"f8c287e8",
  2110 => x"c848bfd4",
  2111 => x"d8f8c280",
  2112 => x"87effe58",
  2113 => x"711e731e",
  2114 => x"9a4a134b",
  2115 => x"7287cb02",
  2116 => x"87e7fe49",
  2117 => x"059a4a13",
  2118 => x"dafe87f5",
  2119 => x"f8c21e87",
  2120 => x"c249bfd4",
  2121 => x"c148d4f8",
  2122 => x"c0c478a1",
  2123 => x"db03a9b7",
  2124 => x"48d4ff87",
  2125 => x"bfd8f8c2",
  2126 => x"d4f8c278",
  2127 => x"f8c249bf",
  2128 => x"a1c148d4",
  2129 => x"b7c0c478",
  2130 => x"87e504a9",
  2131 => x"c848d0ff",
  2132 => x"e0f8c278",
  2133 => x"2678c048",
  2134 => x"0000004f",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00005f5f",
  2138 => x"03030000",
  2139 => x"00030300",
  2140 => x"7f7f1400",
  2141 => x"147f7f14",
  2142 => x"2e240000",
  2143 => x"123a6b6b",
  2144 => x"366a4c00",
  2145 => x"32566c18",
  2146 => x"4f7e3000",
  2147 => x"683a7759",
  2148 => x"04000040",
  2149 => x"00000307",
  2150 => x"1c000000",
  2151 => x"0041633e",
  2152 => x"41000000",
  2153 => x"001c3e63",
  2154 => x"3e2a0800",
  2155 => x"2a3e1c1c",
  2156 => x"08080008",
  2157 => x"08083e3e",
  2158 => x"80000000",
  2159 => x"000060e0",
  2160 => x"08080000",
  2161 => x"08080808",
  2162 => x"00000000",
  2163 => x"00006060",
  2164 => x"30604000",
  2165 => x"03060c18",
  2166 => x"7f3e0001",
  2167 => x"3e7f4d59",
  2168 => x"06040000",
  2169 => x"00007f7f",
  2170 => x"63420000",
  2171 => x"464f5971",
  2172 => x"63220000",
  2173 => x"367f4949",
  2174 => x"161c1800",
  2175 => x"107f7f13",
  2176 => x"67270000",
  2177 => x"397d4545",
  2178 => x"7e3c0000",
  2179 => x"3079494b",
  2180 => x"01010000",
  2181 => x"070f7971",
  2182 => x"7f360000",
  2183 => x"367f4949",
  2184 => x"4f060000",
  2185 => x"1e3f6949",
  2186 => x"00000000",
  2187 => x"00006666",
  2188 => x"80000000",
  2189 => x"000066e6",
  2190 => x"08080000",
  2191 => x"22221414",
  2192 => x"14140000",
  2193 => x"14141414",
  2194 => x"22220000",
  2195 => x"08081414",
  2196 => x"03020000",
  2197 => x"060f5951",
  2198 => x"417f3e00",
  2199 => x"1e1f555d",
  2200 => x"7f7e0000",
  2201 => x"7e7f0909",
  2202 => x"7f7f0000",
  2203 => x"367f4949",
  2204 => x"3e1c0000",
  2205 => x"41414163",
  2206 => x"7f7f0000",
  2207 => x"1c3e6341",
  2208 => x"7f7f0000",
  2209 => x"41414949",
  2210 => x"7f7f0000",
  2211 => x"01010909",
  2212 => x"7f3e0000",
  2213 => x"7a7b4941",
  2214 => x"7f7f0000",
  2215 => x"7f7f0808",
  2216 => x"41000000",
  2217 => x"00417f7f",
  2218 => x"60200000",
  2219 => x"3f7f4040",
  2220 => x"087f7f00",
  2221 => x"4163361c",
  2222 => x"7f7f0000",
  2223 => x"40404040",
  2224 => x"067f7f00",
  2225 => x"7f7f060c",
  2226 => x"067f7f00",
  2227 => x"7f7f180c",
  2228 => x"7f3e0000",
  2229 => x"3e7f4141",
  2230 => x"7f7f0000",
  2231 => x"060f0909",
  2232 => x"417f3e00",
  2233 => x"407e7f61",
  2234 => x"7f7f0000",
  2235 => x"667f1909",
  2236 => x"6f260000",
  2237 => x"327b594d",
  2238 => x"01010000",
  2239 => x"01017f7f",
  2240 => x"7f3f0000",
  2241 => x"3f7f4040",
  2242 => x"3f0f0000",
  2243 => x"0f3f7070",
  2244 => x"307f7f00",
  2245 => x"7f7f3018",
  2246 => x"36634100",
  2247 => x"63361c1c",
  2248 => x"06030141",
  2249 => x"03067c7c",
  2250 => x"59716101",
  2251 => x"4143474d",
  2252 => x"7f000000",
  2253 => x"0041417f",
  2254 => x"06030100",
  2255 => x"6030180c",
  2256 => x"41000040",
  2257 => x"007f7f41",
  2258 => x"060c0800",
  2259 => x"080c0603",
  2260 => x"80808000",
  2261 => x"80808080",
  2262 => x"00000000",
  2263 => x"00040703",
  2264 => x"74200000",
  2265 => x"787c5454",
  2266 => x"7f7f0000",
  2267 => x"387c4444",
  2268 => x"7c380000",
  2269 => x"00444444",
  2270 => x"7c380000",
  2271 => x"7f7f4444",
  2272 => x"7c380000",
  2273 => x"185c5454",
  2274 => x"7e040000",
  2275 => x"0005057f",
  2276 => x"bc180000",
  2277 => x"7cfca4a4",
  2278 => x"7f7f0000",
  2279 => x"787c0404",
  2280 => x"00000000",
  2281 => x"00407d3d",
  2282 => x"80800000",
  2283 => x"007dfd80",
  2284 => x"7f7f0000",
  2285 => x"446c3810",
  2286 => x"00000000",
  2287 => x"00407f3f",
  2288 => x"0c7c7c00",
  2289 => x"787c0c18",
  2290 => x"7c7c0000",
  2291 => x"787c0404",
  2292 => x"7c380000",
  2293 => x"387c4444",
  2294 => x"fcfc0000",
  2295 => x"183c2424",
  2296 => x"3c180000",
  2297 => x"fcfc2424",
  2298 => x"7c7c0000",
  2299 => x"080c0404",
  2300 => x"5c480000",
  2301 => x"20745454",
  2302 => x"3f040000",
  2303 => x"0044447f",
  2304 => x"7c3c0000",
  2305 => x"7c7c4040",
  2306 => x"3c1c0000",
  2307 => x"1c3c6060",
  2308 => x"607c3c00",
  2309 => x"3c7c6030",
  2310 => x"386c4400",
  2311 => x"446c3810",
  2312 => x"bc1c0000",
  2313 => x"1c3c60e0",
  2314 => x"64440000",
  2315 => x"444c5c74",
  2316 => x"08080000",
  2317 => x"4141773e",
  2318 => x"00000000",
  2319 => x"00007f7f",
  2320 => x"41410000",
  2321 => x"08083e77",
  2322 => x"01010200",
  2323 => x"01020203",
  2324 => x"7f7f7f00",
  2325 => x"7f7f7f7f",
  2326 => x"1c080800",
  2327 => x"7f3e3e1c",
  2328 => x"3e7f7f7f",
  2329 => x"081c1c3e",
  2330 => x"18100008",
  2331 => x"10187c7c",
  2332 => x"30100000",
  2333 => x"10307c7c",
  2334 => x"60301000",
  2335 => x"061e7860",
  2336 => x"3c664200",
  2337 => x"42663c18",
  2338 => x"6a387800",
  2339 => x"386cc6c2",
  2340 => x"00006000",
  2341 => x"60000060",
  2342 => x"5b5e0e00",
  2343 => x"1e0e5d5c",
  2344 => x"f8c24c71",
  2345 => x"c04dbff1",
  2346 => x"741ec04b",
  2347 => x"87c702ab",
  2348 => x"c048a6c4",
  2349 => x"c487c578",
  2350 => x"78c148a6",
  2351 => x"731e66c4",
  2352 => x"87dfee49",
  2353 => x"e0c086c8",
  2354 => x"87efef49",
  2355 => x"6a4aa5c4",
  2356 => x"87f0f049",
  2357 => x"cb87c6f1",
  2358 => x"c883c185",
  2359 => x"ff04abb7",
  2360 => x"262687c7",
  2361 => x"264c264d",
  2362 => x"1e4f264b",
  2363 => x"f8c24a71",
  2364 => x"f8c25af5",
  2365 => x"78c748f5",
  2366 => x"87ddfe49",
  2367 => x"731e4f26",
  2368 => x"c04a711e",
  2369 => x"d303aab7",
  2370 => x"dee1c287",
  2371 => x"87c405bf",
  2372 => x"87c24bc1",
  2373 => x"e1c24bc0",
  2374 => x"87c45be2",
  2375 => x"5ae2e1c2",
  2376 => x"bfdee1c2",
  2377 => x"c19ac14a",
  2378 => x"ec49a2c0",
  2379 => x"48fc87e8",
  2380 => x"bfdee1c2",
  2381 => x"87effe78",
  2382 => x"c44a711e",
  2383 => x"49721e66",
  2384 => x"87d2dfff",
  2385 => x"1e4f2626",
  2386 => x"bfdee1c2",
  2387 => x"e5dbff49",
  2388 => x"e9f8c287",
  2389 => x"78bfe848",
  2390 => x"48e5f8c2",
  2391 => x"c278bfec",
  2392 => x"4abfe9f8",
  2393 => x"99ffc349",
  2394 => x"722ab7c8",
  2395 => x"c2b07148",
  2396 => x"2658f1f8",
  2397 => x"5b5e0e4f",
  2398 => x"710e5d5c",
  2399 => x"87c7ff4b",
  2400 => x"48e4f8c2",
  2401 => x"497350c0",
  2402 => x"87cadbff",
  2403 => x"c24c4970",
  2404 => x"49eecb9c",
  2405 => x"7087cfcb",
  2406 => x"f8c24d49",
  2407 => x"05bf97e4",
  2408 => x"d087e4c1",
  2409 => x"f8c24966",
  2410 => x"0599bfed",
  2411 => x"66d487d7",
  2412 => x"e5f8c249",
  2413 => x"cc0599bf",
  2414 => x"ff497387",
  2415 => x"7087d7da",
  2416 => x"c2c10298",
  2417 => x"fd4cc187",
  2418 => x"497587fd",
  2419 => x"7087e3ca",
  2420 => x"87c60298",
  2421 => x"48e4f8c2",
  2422 => x"f8c250c1",
  2423 => x"05bf97e4",
  2424 => x"c287e4c0",
  2425 => x"49bfedf8",
  2426 => x"059966d0",
  2427 => x"c287d6ff",
  2428 => x"49bfe5f8",
  2429 => x"059966d4",
  2430 => x"7387caff",
  2431 => x"d5d9ff49",
  2432 => x"05987087",
  2433 => x"7487fefe",
  2434 => x"87d7fb48",
  2435 => x"5c5b5e0e",
  2436 => x"86f40e5d",
  2437 => x"ec4c4dc0",
  2438 => x"a6c47ebf",
  2439 => x"f1f8c248",
  2440 => x"1ec178bf",
  2441 => x"49c71ec0",
  2442 => x"c887cafd",
  2443 => x"02987086",
  2444 => x"49ff87ce",
  2445 => x"c187c7fb",
  2446 => x"d8ff49da",
  2447 => x"4dc187d8",
  2448 => x"97e4f8c2",
  2449 => x"87c302bf",
  2450 => x"c287c0c9",
  2451 => x"4bbfe9f8",
  2452 => x"bfdee1c2",
  2453 => x"87ebc005",
  2454 => x"ff49fdc3",
  2455 => x"c387f7d7",
  2456 => x"d7ff49fa",
  2457 => x"497387f0",
  2458 => x"7199ffc3",
  2459 => x"fb49c01e",
  2460 => x"497387c6",
  2461 => x"7129b7c8",
  2462 => x"fa49c11e",
  2463 => x"86c887fa",
  2464 => x"c287c1c6",
  2465 => x"4bbfedf8",
  2466 => x"87dd029b",
  2467 => x"bfdae1c2",
  2468 => x"87dec749",
  2469 => x"c4059870",
  2470 => x"d24bc087",
  2471 => x"49e0c287",
  2472 => x"c287c3c7",
  2473 => x"c658dee1",
  2474 => x"dae1c287",
  2475 => x"7378c048",
  2476 => x"0599c249",
  2477 => x"ebc387ce",
  2478 => x"d9d6ff49",
  2479 => x"c2497087",
  2480 => x"87c20299",
  2481 => x"49734cfb",
  2482 => x"ce0599c1",
  2483 => x"49f4c387",
  2484 => x"87c2d6ff",
  2485 => x"99c24970",
  2486 => x"fa87c202",
  2487 => x"c849734c",
  2488 => x"87ce0599",
  2489 => x"ff49f5c3",
  2490 => x"7087ebd5",
  2491 => x"0299c249",
  2492 => x"f8c287d5",
  2493 => x"ca02bff5",
  2494 => x"88c14887",
  2495 => x"58f9f8c2",
  2496 => x"ff87c2c0",
  2497 => x"734dc14c",
  2498 => x"0599c449",
  2499 => x"f2c387ce",
  2500 => x"c1d5ff49",
  2501 => x"c2497087",
  2502 => x"87dc0299",
  2503 => x"bff5f8c2",
  2504 => x"b7c7487e",
  2505 => x"cbc003a8",
  2506 => x"c1486e87",
  2507 => x"f9f8c280",
  2508 => x"87c2c058",
  2509 => x"4dc14cfe",
  2510 => x"ff49fdc3",
  2511 => x"7087d7d4",
  2512 => x"0299c249",
  2513 => x"c287d5c0",
  2514 => x"02bff5f8",
  2515 => x"c287c9c0",
  2516 => x"c048f5f8",
  2517 => x"87c2c078",
  2518 => x"4dc14cfd",
  2519 => x"ff49fac3",
  2520 => x"7087f3d3",
  2521 => x"0299c249",
  2522 => x"c287d9c0",
  2523 => x"48bff5f8",
  2524 => x"03a8b7c7",
  2525 => x"c287c9c0",
  2526 => x"c748f5f8",
  2527 => x"87c2c078",
  2528 => x"4dc14cfc",
  2529 => x"03acb7c0",
  2530 => x"c487d1c0",
  2531 => x"d8c14a66",
  2532 => x"c0026a82",
  2533 => x"4b6a87c6",
  2534 => x"0f734974",
  2535 => x"f0c31ec0",
  2536 => x"49dac11e",
  2537 => x"c887cef7",
  2538 => x"02987086",
  2539 => x"c887e2c0",
  2540 => x"f8c248a6",
  2541 => x"c878bff5",
  2542 => x"91cb4966",
  2543 => x"714866c4",
  2544 => x"6e7e7080",
  2545 => x"c8c002bf",
  2546 => x"4bbf6e87",
  2547 => x"734966c8",
  2548 => x"029d750f",
  2549 => x"c287c8c0",
  2550 => x"49bff5f8",
  2551 => x"c287faf2",
  2552 => x"02bfe2e1",
  2553 => x"4987ddc0",
  2554 => x"7087c7c2",
  2555 => x"d3c00298",
  2556 => x"f5f8c287",
  2557 => x"e0f249bf",
  2558 => x"f449c087",
  2559 => x"e1c287c0",
  2560 => x"78c048e2",
  2561 => x"daf38ef4",
  2562 => x"5b5e0e87",
  2563 => x"1e0e5d5c",
  2564 => x"f8c24c71",
  2565 => x"c149bff1",
  2566 => x"c14da1cd",
  2567 => x"7e6981d1",
  2568 => x"cf029c74",
  2569 => x"4ba5c487",
  2570 => x"f8c27b74",
  2571 => x"f249bff1",
  2572 => x"7b6e87f9",
  2573 => x"c4059c74",
  2574 => x"c24bc087",
  2575 => x"734bc187",
  2576 => x"87faf249",
  2577 => x"c70266d4",
  2578 => x"87da4987",
  2579 => x"87c24a70",
  2580 => x"e1c24ac0",
  2581 => x"f2265ae6",
  2582 => x"000087c9",
  2583 => x"00000000",
  2584 => x"00000000",
  2585 => x"711e0000",
  2586 => x"bfc8ff4a",
  2587 => x"48a17249",
  2588 => x"ff1e4f26",
  2589 => x"fe89bfc8",
  2590 => x"c0c0c0c0",
  2591 => x"c401a9c0",
  2592 => x"c24ac087",
  2593 => x"724ac187",
  2594 => x"1e4f2648",
  2595 => x"bfd9e3c2",
  2596 => x"c2b9c149",
  2597 => x"ff59dde3",
  2598 => x"ffc348d4",
  2599 => x"48d0ff78",
  2600 => x"ff78e1c0",
  2601 => x"78c148d4",
  2602 => x"787131c4",
  2603 => x"c048d0ff",
  2604 => x"4f2678e0",
  2605 => x"cde3c21e",
  2606 => x"d8f3c21e",
  2607 => x"d1fbfd49",
  2608 => x"7086c487",
  2609 => x"87c30298",
  2610 => x"2687c0ff",
  2611 => x"4b35314f",
  2612 => x"20205a48",
  2613 => x"47464320",
  2614 => x"00000000",
  2615 => x"5b5e0e00",
  2616 => x"c20e5d5c",
  2617 => x"4abfe5f8",
  2618 => x"bfc6e5c2",
  2619 => x"bc724c49",
  2620 => x"c5ff4d71",
  2621 => x"4bc087f7",
  2622 => x"99d04974",
  2623 => x"87e7c002",
  2624 => x"c848d0ff",
  2625 => x"d4ff78e1",
  2626 => x"7578c548",
  2627 => x"0299d049",
  2628 => x"f0c387c3",
  2629 => x"f4e5c278",
  2630 => x"11817349",
  2631 => x"08d4ff48",
  2632 => x"48d0ff78",
  2633 => x"c178e0c0",
  2634 => x"c8832d2c",
  2635 => x"c7ff04ab",
  2636 => x"f0c4ff87",
  2637 => x"c6e5c287",
  2638 => x"e5f8c248",
  2639 => x"4d2678bf",
  2640 => x"4b264c26",
  2641 => x"00004f26",
  2642 => x"c11e0000",
  2643 => x"de48d0e7",
  2644 => x"dde5c250",
  2645 => x"fad8fe49",
  2646 => x"2648c087",
  2647 => x"4f544a4f",
  2648 => x"55525455",
  2649 => x"4352414e",
  2650 => x"dff21e00",
  2651 => x"87edfd87",
  2652 => x"4f2687f8",
  2653 => x"25261e16",
  2654 => x"3e3d362e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
