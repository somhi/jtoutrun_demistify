
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"1f",x"ea"),
     1 => (x"48",x"d0",x"ff",x"1e"),
     2 => (x"71",x"78",x"c9",x"c8"),
     3 => (x"08",x"d4",x"ff",x"48"),
     4 => (x"1e",x"4f",x"26",x"78"),
     5 => (x"eb",x"49",x"4a",x"71"),
     6 => (x"48",x"d0",x"ff",x"87"),
     7 => (x"4f",x"26",x"78",x"c8"),
     8 => (x"71",x"1e",x"73",x"1e"),
     9 => (x"e0",x"f7",x"c2",x"4b"),
    10 => (x"87",x"c3",x"02",x"bf"),
    11 => (x"ff",x"87",x"eb",x"c2"),
    12 => (x"c9",x"c8",x"48",x"d0"),
    13 => (x"c0",x"49",x"73",x"78"),
    14 => (x"d4",x"ff",x"b1",x"e0"),
    15 => (x"c2",x"78",x"71",x"48"),
    16 => (x"c0",x"48",x"d4",x"f7"),
    17 => (x"02",x"66",x"c8",x"78"),
    18 => (x"ff",x"c3",x"87",x"c5"),
    19 => (x"c0",x"87",x"c2",x"49"),
    20 => (x"dc",x"f7",x"c2",x"49"),
    21 => (x"02",x"66",x"cc",x"59"),
    22 => (x"d5",x"c5",x"87",x"c6"),
    23 => (x"87",x"c4",x"4a",x"d5"),
    24 => (x"4a",x"ff",x"ff",x"cf"),
    25 => (x"5a",x"e0",x"f7",x"c2"),
    26 => (x"48",x"e0",x"f7",x"c2"),
    27 => (x"87",x"c4",x"78",x"c1"),
    28 => (x"4c",x"26",x"4d",x"26"),
    29 => (x"4f",x"26",x"4b",x"26"),
    30 => (x"5c",x"5b",x"5e",x"0e"),
    31 => (x"4a",x"71",x"0e",x"5d"),
    32 => (x"bf",x"dc",x"f7",x"c2"),
    33 => (x"02",x"9a",x"72",x"4c"),
    34 => (x"c8",x"49",x"87",x"cb"),
    35 => (x"d6",x"c0",x"c2",x"91"),
    36 => (x"c4",x"83",x"71",x"4b"),
    37 => (x"d6",x"c4",x"c2",x"87"),
    38 => (x"13",x"4d",x"c0",x"4b"),
    39 => (x"c2",x"99",x"74",x"49"),
    40 => (x"b9",x"bf",x"d8",x"f7"),
    41 => (x"71",x"48",x"d4",x"ff"),
    42 => (x"2c",x"b7",x"c1",x"78"),
    43 => (x"ad",x"b7",x"c8",x"85"),
    44 => (x"c2",x"87",x"e8",x"04"),
    45 => (x"48",x"bf",x"d4",x"f7"),
    46 => (x"f7",x"c2",x"80",x"c8"),
    47 => (x"ef",x"fe",x"58",x"d8"),
    48 => (x"1e",x"73",x"1e",x"87"),
    49 => (x"4a",x"13",x"4b",x"71"),
    50 => (x"87",x"cb",x"02",x"9a"),
    51 => (x"e7",x"fe",x"49",x"72"),
    52 => (x"9a",x"4a",x"13",x"87"),
    53 => (x"fe",x"87",x"f5",x"05"),
    54 => (x"c2",x"1e",x"87",x"da"),
    55 => (x"49",x"bf",x"d4",x"f7"),
    56 => (x"48",x"d4",x"f7",x"c2"),
    57 => (x"c4",x"78",x"a1",x"c1"),
    58 => (x"03",x"a9",x"b7",x"c0"),
    59 => (x"d4",x"ff",x"87",x"db"),
    60 => (x"d8",x"f7",x"c2",x"48"),
    61 => (x"f7",x"c2",x"78",x"bf"),
    62 => (x"c2",x"49",x"bf",x"d4"),
    63 => (x"c1",x"48",x"d4",x"f7"),
    64 => (x"c0",x"c4",x"78",x"a1"),
    65 => (x"e5",x"04",x"a9",x"b7"),
    66 => (x"48",x"d0",x"ff",x"87"),
    67 => (x"f7",x"c2",x"78",x"c8"),
    68 => (x"78",x"c0",x"48",x"e0"),
    69 => (x"00",x"00",x"4f",x"26"),
    70 => (x"00",x"00",x"00",x"00"),
    71 => (x"00",x"00",x"00",x"00"),
    72 => (x"00",x"5f",x"5f",x"00"),
    73 => (x"03",x"00",x"00",x"00"),
    74 => (x"03",x"03",x"00",x"03"),
    75 => (x"7f",x"14",x"00",x"00"),
    76 => (x"7f",x"7f",x"14",x"7f"),
    77 => (x"24",x"00",x"00",x"14"),
    78 => (x"3a",x"6b",x"6b",x"2e"),
    79 => (x"6a",x"4c",x"00",x"12"),
    80 => (x"56",x"6c",x"18",x"36"),
    81 => (x"7e",x"30",x"00",x"32"),
    82 => (x"3a",x"77",x"59",x"4f"),
    83 => (x"00",x"00",x"40",x"68"),
    84 => (x"00",x"03",x"07",x"04"),
    85 => (x"00",x"00",x"00",x"00"),
    86 => (x"41",x"63",x"3e",x"1c"),
    87 => (x"00",x"00",x"00",x"00"),
    88 => (x"1c",x"3e",x"63",x"41"),
    89 => (x"2a",x"08",x"00",x"00"),
    90 => (x"3e",x"1c",x"1c",x"3e"),
    91 => (x"08",x"00",x"08",x"2a"),
    92 => (x"08",x"3e",x"3e",x"08"),
    93 => (x"00",x"00",x"00",x"08"),
    94 => (x"00",x"60",x"e0",x"80"),
    95 => (x"08",x"00",x"00",x"00"),
    96 => (x"08",x"08",x"08",x"08"),
    97 => (x"00",x"00",x"00",x"08"),
    98 => (x"00",x"60",x"60",x"00"),
    99 => (x"60",x"40",x"00",x"00"),
   100 => (x"06",x"0c",x"18",x"30"),
   101 => (x"3e",x"00",x"01",x"03"),
   102 => (x"7f",x"4d",x"59",x"7f"),
   103 => (x"04",x"00",x"00",x"3e"),
   104 => (x"00",x"7f",x"7f",x"06"),
   105 => (x"42",x"00",x"00",x"00"),
   106 => (x"4f",x"59",x"71",x"63"),
   107 => (x"22",x"00",x"00",x"46"),
   108 => (x"7f",x"49",x"49",x"63"),
   109 => (x"1c",x"18",x"00",x"36"),
   110 => (x"7f",x"7f",x"13",x"16"),
   111 => (x"27",x"00",x"00",x"10"),
   112 => (x"7d",x"45",x"45",x"67"),
   113 => (x"3c",x"00",x"00",x"39"),
   114 => (x"79",x"49",x"4b",x"7e"),
   115 => (x"01",x"00",x"00",x"30"),
   116 => (x"0f",x"79",x"71",x"01"),
   117 => (x"36",x"00",x"00",x"07"),
   118 => (x"7f",x"49",x"49",x"7f"),
   119 => (x"06",x"00",x"00",x"36"),
   120 => (x"3f",x"69",x"49",x"4f"),
   121 => (x"00",x"00",x"00",x"1e"),
   122 => (x"00",x"66",x"66",x"00"),
   123 => (x"00",x"00",x"00",x"00"),
   124 => (x"00",x"66",x"e6",x"80"),
   125 => (x"08",x"00",x"00",x"00"),
   126 => (x"22",x"14",x"14",x"08"),
   127 => (x"14",x"00",x"00",x"22"),
   128 => (x"14",x"14",x"14",x"14"),
   129 => (x"22",x"00",x"00",x"14"),
   130 => (x"08",x"14",x"14",x"22"),
   131 => (x"02",x"00",x"00",x"08"),
   132 => (x"0f",x"59",x"51",x"03"),
   133 => (x"7f",x"3e",x"00",x"06"),
   134 => (x"1f",x"55",x"5d",x"41"),
   135 => (x"7e",x"00",x"00",x"1e"),
   136 => (x"7f",x"09",x"09",x"7f"),
   137 => (x"7f",x"00",x"00",x"7e"),
   138 => (x"7f",x"49",x"49",x"7f"),
   139 => (x"1c",x"00",x"00",x"36"),
   140 => (x"41",x"41",x"63",x"3e"),
   141 => (x"7f",x"00",x"00",x"41"),
   142 => (x"3e",x"63",x"41",x"7f"),
   143 => (x"7f",x"00",x"00",x"1c"),
   144 => (x"41",x"49",x"49",x"7f"),
   145 => (x"7f",x"00",x"00",x"41"),
   146 => (x"01",x"09",x"09",x"7f"),
   147 => (x"3e",x"00",x"00",x"01"),
   148 => (x"7b",x"49",x"41",x"7f"),
   149 => (x"7f",x"00",x"00",x"7a"),
   150 => (x"7f",x"08",x"08",x"7f"),
   151 => (x"00",x"00",x"00",x"7f"),
   152 => (x"41",x"7f",x"7f",x"41"),
   153 => (x"20",x"00",x"00",x"00"),
   154 => (x"7f",x"40",x"40",x"60"),
   155 => (x"7f",x"7f",x"00",x"3f"),
   156 => (x"63",x"36",x"1c",x"08"),
   157 => (x"7f",x"00",x"00",x"41"),
   158 => (x"40",x"40",x"40",x"7f"),
   159 => (x"7f",x"7f",x"00",x"40"),
   160 => (x"7f",x"06",x"0c",x"06"),
   161 => (x"7f",x"7f",x"00",x"7f"),
   162 => (x"7f",x"18",x"0c",x"06"),
   163 => (x"3e",x"00",x"00",x"7f"),
   164 => (x"7f",x"41",x"41",x"7f"),
   165 => (x"7f",x"00",x"00",x"3e"),
   166 => (x"0f",x"09",x"09",x"7f"),
   167 => (x"7f",x"3e",x"00",x"06"),
   168 => (x"7e",x"7f",x"61",x"41"),
   169 => (x"7f",x"00",x"00",x"40"),
   170 => (x"7f",x"19",x"09",x"7f"),
   171 => (x"26",x"00",x"00",x"66"),
   172 => (x"7b",x"59",x"4d",x"6f"),
   173 => (x"01",x"00",x"00",x"32"),
   174 => (x"01",x"7f",x"7f",x"01"),
   175 => (x"3f",x"00",x"00",x"01"),
   176 => (x"7f",x"40",x"40",x"7f"),
   177 => (x"0f",x"00",x"00",x"3f"),
   178 => (x"3f",x"70",x"70",x"3f"),
   179 => (x"7f",x"7f",x"00",x"0f"),
   180 => (x"7f",x"30",x"18",x"30"),
   181 => (x"63",x"41",x"00",x"7f"),
   182 => (x"36",x"1c",x"1c",x"36"),
   183 => (x"03",x"01",x"41",x"63"),
   184 => (x"06",x"7c",x"7c",x"06"),
   185 => (x"71",x"61",x"01",x"03"),
   186 => (x"43",x"47",x"4d",x"59"),
   187 => (x"00",x"00",x"00",x"41"),
   188 => (x"41",x"41",x"7f",x"7f"),
   189 => (x"03",x"01",x"00",x"00"),
   190 => (x"30",x"18",x"0c",x"06"),
   191 => (x"00",x"00",x"40",x"60"),
   192 => (x"7f",x"7f",x"41",x"41"),
   193 => (x"0c",x"08",x"00",x"00"),
   194 => (x"0c",x"06",x"03",x"06"),
   195 => (x"80",x"80",x"00",x"08"),
   196 => (x"80",x"80",x"80",x"80"),
   197 => (x"00",x"00",x"00",x"80"),
   198 => (x"04",x"07",x"03",x"00"),
   199 => (x"20",x"00",x"00",x"00"),
   200 => (x"7c",x"54",x"54",x"74"),
   201 => (x"7f",x"00",x"00",x"78"),
   202 => (x"7c",x"44",x"44",x"7f"),
   203 => (x"38",x"00",x"00",x"38"),
   204 => (x"44",x"44",x"44",x"7c"),
   205 => (x"38",x"00",x"00",x"00"),
   206 => (x"7f",x"44",x"44",x"7c"),
   207 => (x"38",x"00",x"00",x"7f"),
   208 => (x"5c",x"54",x"54",x"7c"),
   209 => (x"04",x"00",x"00",x"18"),
   210 => (x"05",x"05",x"7f",x"7e"),
   211 => (x"18",x"00",x"00",x"00"),
   212 => (x"fc",x"a4",x"a4",x"bc"),
   213 => (x"7f",x"00",x"00",x"7c"),
   214 => (x"7c",x"04",x"04",x"7f"),
   215 => (x"00",x"00",x"00",x"78"),
   216 => (x"40",x"7d",x"3d",x"00"),
   217 => (x"80",x"00",x"00",x"00"),
   218 => (x"7d",x"fd",x"80",x"80"),
   219 => (x"7f",x"00",x"00",x"00"),
   220 => (x"6c",x"38",x"10",x"7f"),
   221 => (x"00",x"00",x"00",x"44"),
   222 => (x"40",x"7f",x"3f",x"00"),
   223 => (x"7c",x"7c",x"00",x"00"),
   224 => (x"7c",x"0c",x"18",x"0c"),
   225 => (x"7c",x"00",x"00",x"78"),
   226 => (x"7c",x"04",x"04",x"7c"),
   227 => (x"38",x"00",x"00",x"78"),
   228 => (x"7c",x"44",x"44",x"7c"),
   229 => (x"fc",x"00",x"00",x"38"),
   230 => (x"3c",x"24",x"24",x"fc"),
   231 => (x"18",x"00",x"00",x"18"),
   232 => (x"fc",x"24",x"24",x"3c"),
   233 => (x"7c",x"00",x"00",x"fc"),
   234 => (x"0c",x"04",x"04",x"7c"),
   235 => (x"48",x"00",x"00",x"08"),
   236 => (x"74",x"54",x"54",x"5c"),
   237 => (x"04",x"00",x"00",x"20"),
   238 => (x"44",x"44",x"7f",x"3f"),
   239 => (x"3c",x"00",x"00",x"00"),
   240 => (x"7c",x"40",x"40",x"7c"),
   241 => (x"1c",x"00",x"00",x"7c"),
   242 => (x"3c",x"60",x"60",x"3c"),
   243 => (x"7c",x"3c",x"00",x"1c"),
   244 => (x"7c",x"60",x"30",x"60"),
   245 => (x"6c",x"44",x"00",x"3c"),
   246 => (x"6c",x"38",x"10",x"38"),
   247 => (x"1c",x"00",x"00",x"44"),
   248 => (x"3c",x"60",x"e0",x"bc"),
   249 => (x"44",x"00",x"00",x"1c"),
   250 => (x"4c",x"5c",x"74",x"64"),
   251 => (x"08",x"00",x"00",x"44"),
   252 => (x"41",x"77",x"3e",x"08"),
   253 => (x"00",x"00",x"00",x"41"),
   254 => (x"00",x"7f",x"7f",x"00"),
   255 => (x"41",x"00",x"00",x"00"),
   256 => (x"08",x"3e",x"77",x"41"),
   257 => (x"01",x"02",x"00",x"08"),
   258 => (x"02",x"02",x"03",x"01"),
   259 => (x"7f",x"7f",x"00",x"01"),
   260 => (x"7f",x"7f",x"7f",x"7f"),
   261 => (x"08",x"08",x"00",x"7f"),
   262 => (x"3e",x"3e",x"1c",x"1c"),
   263 => (x"7f",x"7f",x"7f",x"7f"),
   264 => (x"1c",x"1c",x"3e",x"3e"),
   265 => (x"10",x"00",x"08",x"08"),
   266 => (x"18",x"7c",x"7c",x"18"),
   267 => (x"10",x"00",x"00",x"10"),
   268 => (x"30",x"7c",x"7c",x"30"),
   269 => (x"30",x"10",x"00",x"10"),
   270 => (x"1e",x"78",x"60",x"60"),
   271 => (x"66",x"42",x"00",x"06"),
   272 => (x"66",x"3c",x"18",x"3c"),
   273 => (x"38",x"78",x"00",x"42"),
   274 => (x"6c",x"c6",x"c2",x"6a"),
   275 => (x"00",x"60",x"00",x"38"),
   276 => (x"00",x"00",x"60",x"00"),
   277 => (x"5e",x"0e",x"00",x"60"),
   278 => (x"0e",x"5d",x"5c",x"5b"),
   279 => (x"c2",x"4c",x"71",x"1e"),
   280 => (x"4d",x"bf",x"f1",x"f7"),
   281 => (x"1e",x"c0",x"4b",x"c0"),
   282 => (x"c7",x"02",x"ab",x"74"),
   283 => (x"48",x"a6",x"c4",x"87"),
   284 => (x"87",x"c5",x"78",x"c0"),
   285 => (x"c1",x"48",x"a6",x"c4"),
   286 => (x"1e",x"66",x"c4",x"78"),
   287 => (x"df",x"ee",x"49",x"73"),
   288 => (x"c0",x"86",x"c8",x"87"),
   289 => (x"ef",x"ef",x"49",x"e0"),
   290 => (x"4a",x"a5",x"c4",x"87"),
   291 => (x"f0",x"f0",x"49",x"6a"),
   292 => (x"87",x"c6",x"f1",x"87"),
   293 => (x"83",x"c1",x"85",x"cb"),
   294 => (x"04",x"ab",x"b7",x"c8"),
   295 => (x"26",x"87",x"c7",x"ff"),
   296 => (x"4c",x"26",x"4d",x"26"),
   297 => (x"4f",x"26",x"4b",x"26"),
   298 => (x"c2",x"4a",x"71",x"1e"),
   299 => (x"c2",x"5a",x"f5",x"f7"),
   300 => (x"c7",x"48",x"f5",x"f7"),
   301 => (x"dd",x"fe",x"49",x"78"),
   302 => (x"1e",x"4f",x"26",x"87"),
   303 => (x"4a",x"71",x"1e",x"73"),
   304 => (x"03",x"aa",x"b7",x"c0"),
   305 => (x"e0",x"c2",x"87",x"d3"),
   306 => (x"c4",x"05",x"bf",x"db"),
   307 => (x"c2",x"4b",x"c1",x"87"),
   308 => (x"c2",x"4b",x"c0",x"87"),
   309 => (x"c4",x"5b",x"df",x"e0"),
   310 => (x"df",x"e0",x"c2",x"87"),
   311 => (x"db",x"e0",x"c2",x"5a"),
   312 => (x"9a",x"c1",x"4a",x"bf"),
   313 => (x"49",x"a2",x"c0",x"c1"),
   314 => (x"fc",x"87",x"e8",x"ec"),
   315 => (x"db",x"e0",x"c2",x"48"),
   316 => (x"ef",x"fe",x"78",x"bf"),
   317 => (x"4a",x"71",x"1e",x"87"),
   318 => (x"72",x"1e",x"66",x"c4"),
   319 => (x"e9",x"df",x"ff",x"49"),
   320 => (x"4f",x"26",x"26",x"87"),
   321 => (x"db",x"e0",x"c2",x"1e"),
   322 => (x"dc",x"ff",x"49",x"bf"),
   323 => (x"f7",x"c2",x"87",x"d9"),
   324 => (x"bf",x"e8",x"48",x"e9"),
   325 => (x"e5",x"f7",x"c2",x"78"),
   326 => (x"78",x"bf",x"ec",x"48"),
   327 => (x"bf",x"e9",x"f7",x"c2"),
   328 => (x"ff",x"c3",x"49",x"4a"),
   329 => (x"2a",x"b7",x"c8",x"99"),
   330 => (x"b0",x"71",x"48",x"72"),
   331 => (x"58",x"f1",x"f7",x"c2"),
   332 => (x"5e",x"0e",x"4f",x"26"),
   333 => (x"0e",x"5d",x"5c",x"5b"),
   334 => (x"c7",x"ff",x"4b",x"71"),
   335 => (x"e4",x"f7",x"c2",x"87"),
   336 => (x"73",x"50",x"c0",x"48"),
   337 => (x"fe",x"db",x"ff",x"49"),
   338 => (x"4c",x"49",x"70",x"87"),
   339 => (x"ee",x"cb",x"9c",x"c2"),
   340 => (x"87",x"cf",x"cb",x"49"),
   341 => (x"c2",x"4d",x"49",x"70"),
   342 => (x"bf",x"97",x"e4",x"f7"),
   343 => (x"87",x"e4",x"c1",x"05"),
   344 => (x"c2",x"49",x"66",x"d0"),
   345 => (x"99",x"bf",x"ed",x"f7"),
   346 => (x"d4",x"87",x"d7",x"05"),
   347 => (x"f7",x"c2",x"49",x"66"),
   348 => (x"05",x"99",x"bf",x"e5"),
   349 => (x"49",x"73",x"87",x"cc"),
   350 => (x"87",x"cb",x"db",x"ff"),
   351 => (x"c1",x"02",x"98",x"70"),
   352 => (x"4c",x"c1",x"87",x"c2"),
   353 => (x"75",x"87",x"fd",x"fd"),
   354 => (x"87",x"e3",x"ca",x"49"),
   355 => (x"c6",x"02",x"98",x"70"),
   356 => (x"e4",x"f7",x"c2",x"87"),
   357 => (x"c2",x"50",x"c1",x"48"),
   358 => (x"bf",x"97",x"e4",x"f7"),
   359 => (x"87",x"e4",x"c0",x"05"),
   360 => (x"bf",x"ed",x"f7",x"c2"),
   361 => (x"99",x"66",x"d0",x"49"),
   362 => (x"87",x"d6",x"ff",x"05"),
   363 => (x"bf",x"e5",x"f7",x"c2"),
   364 => (x"99",x"66",x"d4",x"49"),
   365 => (x"87",x"ca",x"ff",x"05"),
   366 => (x"da",x"ff",x"49",x"73"),
   367 => (x"98",x"70",x"87",x"c9"),
   368 => (x"87",x"fe",x"fe",x"05"),
   369 => (x"d7",x"fb",x"48",x"74"),
   370 => (x"5b",x"5e",x"0e",x"87"),
   371 => (x"f4",x"0e",x"5d",x"5c"),
   372 => (x"4c",x"4d",x"c0",x"86"),
   373 => (x"c4",x"7e",x"bf",x"ec"),
   374 => (x"f7",x"c2",x"48",x"a6"),
   375 => (x"c1",x"78",x"bf",x"f1"),
   376 => (x"c7",x"1e",x"c0",x"1e"),
   377 => (x"87",x"ca",x"fd",x"49"),
   378 => (x"98",x"70",x"86",x"c8"),
   379 => (x"ff",x"87",x"ce",x"02"),
   380 => (x"87",x"c7",x"fb",x"49"),
   381 => (x"ff",x"49",x"da",x"c1"),
   382 => (x"c1",x"87",x"cc",x"d9"),
   383 => (x"e4",x"f7",x"c2",x"4d"),
   384 => (x"c3",x"02",x"bf",x"97"),
   385 => (x"87",x"c0",x"c9",x"87"),
   386 => (x"bf",x"e9",x"f7",x"c2"),
   387 => (x"db",x"e0",x"c2",x"4b"),
   388 => (x"eb",x"c0",x"05",x"bf"),
   389 => (x"49",x"fd",x"c3",x"87"),
   390 => (x"87",x"eb",x"d8",x"ff"),
   391 => (x"ff",x"49",x"fa",x"c3"),
   392 => (x"73",x"87",x"e4",x"d8"),
   393 => (x"99",x"ff",x"c3",x"49"),
   394 => (x"49",x"c0",x"1e",x"71"),
   395 => (x"73",x"87",x"c6",x"fb"),
   396 => (x"29",x"b7",x"c8",x"49"),
   397 => (x"49",x"c1",x"1e",x"71"),
   398 => (x"c8",x"87",x"fa",x"fa"),
   399 => (x"87",x"c1",x"c6",x"86"),
   400 => (x"bf",x"ed",x"f7",x"c2"),
   401 => (x"dd",x"02",x"9b",x"4b"),
   402 => (x"d7",x"e0",x"c2",x"87"),
   403 => (x"de",x"c7",x"49",x"bf"),
   404 => (x"05",x"98",x"70",x"87"),
   405 => (x"4b",x"c0",x"87",x"c4"),
   406 => (x"e0",x"c2",x"87",x"d2"),
   407 => (x"87",x"c3",x"c7",x"49"),
   408 => (x"58",x"db",x"e0",x"c2"),
   409 => (x"e0",x"c2",x"87",x"c6"),
   410 => (x"78",x"c0",x"48",x"d7"),
   411 => (x"99",x"c2",x"49",x"73"),
   412 => (x"c3",x"87",x"ce",x"05"),
   413 => (x"d7",x"ff",x"49",x"eb"),
   414 => (x"49",x"70",x"87",x"cd"),
   415 => (x"c2",x"02",x"99",x"c2"),
   416 => (x"73",x"4c",x"fb",x"87"),
   417 => (x"05",x"99",x"c1",x"49"),
   418 => (x"f4",x"c3",x"87",x"ce"),
   419 => (x"f6",x"d6",x"ff",x"49"),
   420 => (x"c2",x"49",x"70",x"87"),
   421 => (x"87",x"c2",x"02",x"99"),
   422 => (x"49",x"73",x"4c",x"fa"),
   423 => (x"ce",x"05",x"99",x"c8"),
   424 => (x"49",x"f5",x"c3",x"87"),
   425 => (x"87",x"df",x"d6",x"ff"),
   426 => (x"99",x"c2",x"49",x"70"),
   427 => (x"c2",x"87",x"d5",x"02"),
   428 => (x"02",x"bf",x"f5",x"f7"),
   429 => (x"c1",x"48",x"87",x"ca"),
   430 => (x"f9",x"f7",x"c2",x"88"),
   431 => (x"87",x"c2",x"c0",x"58"),
   432 => (x"4d",x"c1",x"4c",x"ff"),
   433 => (x"99",x"c4",x"49",x"73"),
   434 => (x"c3",x"87",x"ce",x"05"),
   435 => (x"d5",x"ff",x"49",x"f2"),
   436 => (x"49",x"70",x"87",x"f5"),
   437 => (x"dc",x"02",x"99",x"c2"),
   438 => (x"f5",x"f7",x"c2",x"87"),
   439 => (x"c7",x"48",x"7e",x"bf"),
   440 => (x"c0",x"03",x"a8",x"b7"),
   441 => (x"48",x"6e",x"87",x"cb"),
   442 => (x"f7",x"c2",x"80",x"c1"),
   443 => (x"c2",x"c0",x"58",x"f9"),
   444 => (x"c1",x"4c",x"fe",x"87"),
   445 => (x"49",x"fd",x"c3",x"4d"),
   446 => (x"87",x"cb",x"d5",x"ff"),
   447 => (x"99",x"c2",x"49",x"70"),
   448 => (x"87",x"d5",x"c0",x"02"),
   449 => (x"bf",x"f5",x"f7",x"c2"),
   450 => (x"87",x"c9",x"c0",x"02"),
   451 => (x"48",x"f5",x"f7",x"c2"),
   452 => (x"c2",x"c0",x"78",x"c0"),
   453 => (x"c1",x"4c",x"fd",x"87"),
   454 => (x"49",x"fa",x"c3",x"4d"),
   455 => (x"87",x"e7",x"d4",x"ff"),
   456 => (x"99",x"c2",x"49",x"70"),
   457 => (x"87",x"d9",x"c0",x"02"),
   458 => (x"bf",x"f5",x"f7",x"c2"),
   459 => (x"a8",x"b7",x"c7",x"48"),
   460 => (x"87",x"c9",x"c0",x"03"),
   461 => (x"48",x"f5",x"f7",x"c2"),
   462 => (x"c2",x"c0",x"78",x"c7"),
   463 => (x"c1",x"4c",x"fc",x"87"),
   464 => (x"ac",x"b7",x"c0",x"4d"),
   465 => (x"87",x"d1",x"c0",x"03"),
   466 => (x"c1",x"4a",x"66",x"c4"),
   467 => (x"02",x"6a",x"82",x"d8"),
   468 => (x"6a",x"87",x"c6",x"c0"),
   469 => (x"73",x"49",x"74",x"4b"),
   470 => (x"c3",x"1e",x"c0",x"0f"),
   471 => (x"da",x"c1",x"1e",x"f0"),
   472 => (x"87",x"ce",x"f7",x"49"),
   473 => (x"98",x"70",x"86",x"c8"),
   474 => (x"87",x"e2",x"c0",x"02"),
   475 => (x"c2",x"48",x"a6",x"c8"),
   476 => (x"78",x"bf",x"f5",x"f7"),
   477 => (x"cb",x"49",x"66",x"c8"),
   478 => (x"48",x"66",x"c4",x"91"),
   479 => (x"7e",x"70",x"80",x"71"),
   480 => (x"c0",x"02",x"bf",x"6e"),
   481 => (x"bf",x"6e",x"87",x"c8"),
   482 => (x"49",x"66",x"c8",x"4b"),
   483 => (x"9d",x"75",x"0f",x"73"),
   484 => (x"87",x"c8",x"c0",x"02"),
   485 => (x"bf",x"f5",x"f7",x"c2"),
   486 => (x"87",x"fa",x"f2",x"49"),
   487 => (x"bf",x"df",x"e0",x"c2"),
   488 => (x"87",x"dd",x"c0",x"02"),
   489 => (x"87",x"c7",x"c2",x"49"),
   490 => (x"c0",x"02",x"98",x"70"),
   491 => (x"f7",x"c2",x"87",x"d3"),
   492 => (x"f2",x"49",x"bf",x"f5"),
   493 => (x"49",x"c0",x"87",x"e0"),
   494 => (x"c2",x"87",x"c0",x"f4"),
   495 => (x"c0",x"48",x"df",x"e0"),
   496 => (x"f3",x"8e",x"f4",x"78"),
   497 => (x"5e",x"0e",x"87",x"da"),
   498 => (x"0e",x"5d",x"5c",x"5b"),
   499 => (x"c2",x"4c",x"71",x"1e"),
   500 => (x"49",x"bf",x"f1",x"f7"),
   501 => (x"4d",x"a1",x"cd",x"c1"),
   502 => (x"69",x"81",x"d1",x"c1"),
   503 => (x"02",x"9c",x"74",x"7e"),
   504 => (x"a5",x"c4",x"87",x"cf"),
   505 => (x"c2",x"7b",x"74",x"4b"),
   506 => (x"49",x"bf",x"f1",x"f7"),
   507 => (x"6e",x"87",x"f9",x"f2"),
   508 => (x"05",x"9c",x"74",x"7b"),
   509 => (x"4b",x"c0",x"87",x"c4"),
   510 => (x"4b",x"c1",x"87",x"c2"),
   511 => (x"fa",x"f2",x"49",x"73"),
   512 => (x"02",x"66",x"d4",x"87"),
   513 => (x"da",x"49",x"87",x"c7"),
   514 => (x"c2",x"4a",x"70",x"87"),
   515 => (x"c2",x"4a",x"c0",x"87"),
   516 => (x"26",x"5a",x"e3",x"e0"),
   517 => (x"00",x"87",x"c9",x"f2"),
   518 => (x"00",x"00",x"00",x"00"),
   519 => (x"00",x"00",x"00",x"00"),
   520 => (x"1e",x"00",x"00",x"00"),
   521 => (x"c8",x"ff",x"4a",x"71"),
   522 => (x"a1",x"72",x"49",x"bf"),
   523 => (x"1e",x"4f",x"26",x"48"),
   524 => (x"89",x"bf",x"c8",x"ff"),
   525 => (x"c0",x"c0",x"c0",x"fe"),
   526 => (x"01",x"a9",x"c0",x"c0"),
   527 => (x"4a",x"c0",x"87",x"c4"),
   528 => (x"4a",x"c1",x"87",x"c2"),
   529 => (x"4f",x"26",x"48",x"72"),
   530 => (x"d6",x"e2",x"c2",x"1e"),
   531 => (x"b9",x"c1",x"49",x"bf"),
   532 => (x"59",x"da",x"e2",x"c2"),
   533 => (x"c3",x"48",x"d4",x"ff"),
   534 => (x"d0",x"ff",x"78",x"ff"),
   535 => (x"78",x"e1",x"c0",x"48"),
   536 => (x"c1",x"48",x"d4",x"ff"),
   537 => (x"71",x"31",x"c4",x"78"),
   538 => (x"48",x"d0",x"ff",x"78"),
   539 => (x"26",x"78",x"e0",x"c0"),
   540 => (x"e2",x"c2",x"1e",x"4f"),
   541 => (x"f2",x"c2",x"1e",x"ca"),
   542 => (x"fc",x"fd",x"49",x"d8"),
   543 => (x"86",x"c4",x"87",x"c7"),
   544 => (x"c3",x"02",x"98",x"70"),
   545 => (x"87",x"c0",x"ff",x"87"),
   546 => (x"35",x"31",x"4f",x"26"),
   547 => (x"20",x"5a",x"48",x"4b"),
   548 => (x"46",x"43",x"20",x"20"),
   549 => (x"00",x"00",x"00",x"47"),
   550 => (x"5e",x"0e",x"00",x"00"),
   551 => (x"0e",x"5d",x"5c",x"5b"),
   552 => (x"bf",x"e5",x"f7",x"c2"),
   553 => (x"c3",x"e4",x"c2",x"4a"),
   554 => (x"72",x"4c",x"49",x"bf"),
   555 => (x"ff",x"4d",x"71",x"bc"),
   556 => (x"c0",x"87",x"eb",x"c6"),
   557 => (x"d0",x"49",x"74",x"4b"),
   558 => (x"e7",x"c0",x"02",x"99"),
   559 => (x"48",x"d0",x"ff",x"87"),
   560 => (x"ff",x"78",x"e1",x"c8"),
   561 => (x"78",x"c5",x"48",x"d4"),
   562 => (x"99",x"d0",x"49",x"75"),
   563 => (x"c3",x"87",x"c3",x"02"),
   564 => (x"e4",x"c2",x"78",x"f0"),
   565 => (x"81",x"73",x"49",x"f1"),
   566 => (x"d4",x"ff",x"48",x"11"),
   567 => (x"d0",x"ff",x"78",x"08"),
   568 => (x"78",x"e0",x"c0",x"48"),
   569 => (x"83",x"2d",x"2c",x"c1"),
   570 => (x"ff",x"04",x"ab",x"c8"),
   571 => (x"c5",x"ff",x"87",x"c7"),
   572 => (x"e4",x"c2",x"87",x"e4"),
   573 => (x"f7",x"c2",x"48",x"c3"),
   574 => (x"26",x"78",x"bf",x"e5"),
   575 => (x"26",x"4c",x"26",x"4d"),
   576 => (x"00",x"4f",x"26",x"4b"),
   577 => (x"1e",x"00",x"00",x"00"),
   578 => (x"48",x"c9",x"e7",x"c1"),
   579 => (x"e4",x"c2",x"50",x"de"),
   580 => (x"d9",x"fe",x"49",x"da"),
   581 => (x"48",x"c0",x"87",x"f1"),
   582 => (x"54",x"4a",x"4f",x"26"),
   583 => (x"52",x"54",x"55",x"4f"),
   584 => (x"52",x"41",x"4e",x"55"),
   585 => (x"f2",x"1e",x"00",x"43"),
   586 => (x"ed",x"fd",x"87",x"df"),
   587 => (x"26",x"87",x"f8",x"87"),
   588 => (x"26",x"1e",x"16",x"4f"),
   589 => (x"3d",x"36",x"2e",x"25"),
   590 => (x"3d",x"36",x"2e",x"3e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

