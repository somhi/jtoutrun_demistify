library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"ed00001f",
     1 => x"1e00001f",
     2 => x"c848d0ff",
     3 => x"487178c9",
     4 => x"7808d4ff",
     5 => x"711e4f26",
     6 => x"87eb494a",
     7 => x"c848d0ff",
     8 => x"1e4f2678",
     9 => x"4b711e73",
    10 => x"bfe0f7c2",
    11 => x"c287c302",
    12 => x"d0ff87eb",
    13 => x"78c9c848",
    14 => x"e0c04973",
    15 => x"48d4ffb1",
    16 => x"f7c27871",
    17 => x"78c048d4",
    18 => x"c50266c8",
    19 => x"49ffc387",
    20 => x"49c087c2",
    21 => x"59dcf7c2",
    22 => x"c60266cc",
    23 => x"d5d5c587",
    24 => x"cf87c44a",
    25 => x"c24affff",
    26 => x"c25ae0f7",
    27 => x"c148e0f7",
    28 => x"2687c478",
    29 => x"264c264d",
    30 => x"0e4f264b",
    31 => x"5d5c5b5e",
    32 => x"c24a710e",
    33 => x"4cbfdcf7",
    34 => x"cb029a72",
    35 => x"91c84987",
    36 => x"4bd9c0c2",
    37 => x"87c48371",
    38 => x"4bd9c4c2",
    39 => x"49134dc0",
    40 => x"f7c29974",
    41 => x"ffb9bfd8",
    42 => x"787148d4",
    43 => x"852cb7c1",
    44 => x"04adb7c8",
    45 => x"f7c287e8",
    46 => x"c848bfd4",
    47 => x"d8f7c280",
    48 => x"87effe58",
    49 => x"711e731e",
    50 => x"9a4a134b",
    51 => x"7287cb02",
    52 => x"87e7fe49",
    53 => x"059a4a13",
    54 => x"dafe87f5",
    55 => x"f7c21e87",
    56 => x"c249bfd4",
    57 => x"c148d4f7",
    58 => x"c0c478a1",
    59 => x"db03a9b7",
    60 => x"48d4ff87",
    61 => x"bfd8f7c2",
    62 => x"d4f7c278",
    63 => x"f7c249bf",
    64 => x"a1c148d4",
    65 => x"b7c0c478",
    66 => x"87e504a9",
    67 => x"c848d0ff",
    68 => x"e0f7c278",
    69 => x"2678c048",
    70 => x"0000004f",
    71 => x"00000000",
    72 => x"00000000",
    73 => x"00005f5f",
    74 => x"03030000",
    75 => x"00030300",
    76 => x"7f7f1400",
    77 => x"147f7f14",
    78 => x"2e240000",
    79 => x"123a6b6b",
    80 => x"366a4c00",
    81 => x"32566c18",
    82 => x"4f7e3000",
    83 => x"683a7759",
    84 => x"04000040",
    85 => x"00000307",
    86 => x"1c000000",
    87 => x"0041633e",
    88 => x"41000000",
    89 => x"001c3e63",
    90 => x"3e2a0800",
    91 => x"2a3e1c1c",
    92 => x"08080008",
    93 => x"08083e3e",
    94 => x"80000000",
    95 => x"000060e0",
    96 => x"08080000",
    97 => x"08080808",
    98 => x"00000000",
    99 => x"00006060",
   100 => x"30604000",
   101 => x"03060c18",
   102 => x"7f3e0001",
   103 => x"3e7f4d59",
   104 => x"06040000",
   105 => x"00007f7f",
   106 => x"63420000",
   107 => x"464f5971",
   108 => x"63220000",
   109 => x"367f4949",
   110 => x"161c1800",
   111 => x"107f7f13",
   112 => x"67270000",
   113 => x"397d4545",
   114 => x"7e3c0000",
   115 => x"3079494b",
   116 => x"01010000",
   117 => x"070f7971",
   118 => x"7f360000",
   119 => x"367f4949",
   120 => x"4f060000",
   121 => x"1e3f6949",
   122 => x"00000000",
   123 => x"00006666",
   124 => x"80000000",
   125 => x"000066e6",
   126 => x"08080000",
   127 => x"22221414",
   128 => x"14140000",
   129 => x"14141414",
   130 => x"22220000",
   131 => x"08081414",
   132 => x"03020000",
   133 => x"060f5951",
   134 => x"417f3e00",
   135 => x"1e1f555d",
   136 => x"7f7e0000",
   137 => x"7e7f0909",
   138 => x"7f7f0000",
   139 => x"367f4949",
   140 => x"3e1c0000",
   141 => x"41414163",
   142 => x"7f7f0000",
   143 => x"1c3e6341",
   144 => x"7f7f0000",
   145 => x"41414949",
   146 => x"7f7f0000",
   147 => x"01010909",
   148 => x"7f3e0000",
   149 => x"7a7b4941",
   150 => x"7f7f0000",
   151 => x"7f7f0808",
   152 => x"41000000",
   153 => x"00417f7f",
   154 => x"60200000",
   155 => x"3f7f4040",
   156 => x"087f7f00",
   157 => x"4163361c",
   158 => x"7f7f0000",
   159 => x"40404040",
   160 => x"067f7f00",
   161 => x"7f7f060c",
   162 => x"067f7f00",
   163 => x"7f7f180c",
   164 => x"7f3e0000",
   165 => x"3e7f4141",
   166 => x"7f7f0000",
   167 => x"060f0909",
   168 => x"417f3e00",
   169 => x"407e7f61",
   170 => x"7f7f0000",
   171 => x"667f1909",
   172 => x"6f260000",
   173 => x"327b594d",
   174 => x"01010000",
   175 => x"01017f7f",
   176 => x"7f3f0000",
   177 => x"3f7f4040",
   178 => x"3f0f0000",
   179 => x"0f3f7070",
   180 => x"307f7f00",
   181 => x"7f7f3018",
   182 => x"36634100",
   183 => x"63361c1c",
   184 => x"06030141",
   185 => x"03067c7c",
   186 => x"59716101",
   187 => x"4143474d",
   188 => x"7f000000",
   189 => x"0041417f",
   190 => x"06030100",
   191 => x"6030180c",
   192 => x"41000040",
   193 => x"007f7f41",
   194 => x"060c0800",
   195 => x"080c0603",
   196 => x"80808000",
   197 => x"80808080",
   198 => x"00000000",
   199 => x"00040703",
   200 => x"74200000",
   201 => x"787c5454",
   202 => x"7f7f0000",
   203 => x"387c4444",
   204 => x"7c380000",
   205 => x"00444444",
   206 => x"7c380000",
   207 => x"7f7f4444",
   208 => x"7c380000",
   209 => x"185c5454",
   210 => x"7e040000",
   211 => x"0005057f",
   212 => x"bc180000",
   213 => x"7cfca4a4",
   214 => x"7f7f0000",
   215 => x"787c0404",
   216 => x"00000000",
   217 => x"00407d3d",
   218 => x"80800000",
   219 => x"007dfd80",
   220 => x"7f7f0000",
   221 => x"446c3810",
   222 => x"00000000",
   223 => x"00407f3f",
   224 => x"0c7c7c00",
   225 => x"787c0c18",
   226 => x"7c7c0000",
   227 => x"787c0404",
   228 => x"7c380000",
   229 => x"387c4444",
   230 => x"fcfc0000",
   231 => x"183c2424",
   232 => x"3c180000",
   233 => x"fcfc2424",
   234 => x"7c7c0000",
   235 => x"080c0404",
   236 => x"5c480000",
   237 => x"20745454",
   238 => x"3f040000",
   239 => x"0044447f",
   240 => x"7c3c0000",
   241 => x"7c7c4040",
   242 => x"3c1c0000",
   243 => x"1c3c6060",
   244 => x"607c3c00",
   245 => x"3c7c6030",
   246 => x"386c4400",
   247 => x"446c3810",
   248 => x"bc1c0000",
   249 => x"1c3c60e0",
   250 => x"64440000",
   251 => x"444c5c74",
   252 => x"08080000",
   253 => x"4141773e",
   254 => x"00000000",
   255 => x"00007f7f",
   256 => x"41410000",
   257 => x"08083e77",
   258 => x"01010200",
   259 => x"01020203",
   260 => x"7f7f7f00",
   261 => x"7f7f7f7f",
   262 => x"1c080800",
   263 => x"7f3e3e1c",
   264 => x"3e7f7f7f",
   265 => x"081c1c3e",
   266 => x"18100008",
   267 => x"10187c7c",
   268 => x"30100000",
   269 => x"10307c7c",
   270 => x"60301000",
   271 => x"061e7860",
   272 => x"3c664200",
   273 => x"42663c18",
   274 => x"6a387800",
   275 => x"386cc6c2",
   276 => x"00006000",
   277 => x"60000060",
   278 => x"5b5e0e00",
   279 => x"1e0e5d5c",
   280 => x"f7c24c71",
   281 => x"c04dbff1",
   282 => x"741ec04b",
   283 => x"87c702ab",
   284 => x"c048a6c4",
   285 => x"c487c578",
   286 => x"78c148a6",
   287 => x"731e66c4",
   288 => x"87dfee49",
   289 => x"e0c086c8",
   290 => x"87efef49",
   291 => x"6a4aa5c4",
   292 => x"87f0f049",
   293 => x"cb87c6f1",
   294 => x"c883c185",
   295 => x"ff04abb7",
   296 => x"262687c7",
   297 => x"264c264d",
   298 => x"1e4f264b",
   299 => x"f7c24a71",
   300 => x"f7c25af5",
   301 => x"78c748f5",
   302 => x"87ddfe49",
   303 => x"731e4f26",
   304 => x"c04a711e",
   305 => x"d303aab7",
   306 => x"dee0c287",
   307 => x"87c405bf",
   308 => x"87c24bc1",
   309 => x"e0c24bc0",
   310 => x"87c45be2",
   311 => x"5ae2e0c2",
   312 => x"bfdee0c2",
   313 => x"c19ac14a",
   314 => x"ec49a2c0",
   315 => x"48fc87e8",
   316 => x"bfdee0c2",
   317 => x"87effe78",
   318 => x"c44a711e",
   319 => x"49721e66",
   320 => x"87e9dfff",
   321 => x"1e4f2626",
   322 => x"bfdee0c2",
   323 => x"d9dcff49",
   324 => x"e9f7c287",
   325 => x"78bfe848",
   326 => x"48e5f7c2",
   327 => x"c278bfec",
   328 => x"4abfe9f7",
   329 => x"99ffc349",
   330 => x"722ab7c8",
   331 => x"c2b07148",
   332 => x"2658f1f7",
   333 => x"5b5e0e4f",
   334 => x"710e5d5c",
   335 => x"87c7ff4b",
   336 => x"48e4f7c2",
   337 => x"497350c0",
   338 => x"87fedbff",
   339 => x"c24c4970",
   340 => x"49eecb9c",
   341 => x"7087cfcb",
   342 => x"f7c24d49",
   343 => x"05bf97e4",
   344 => x"d087e4c1",
   345 => x"f7c24966",
   346 => x"0599bfed",
   347 => x"66d487d7",
   348 => x"e5f7c249",
   349 => x"cc0599bf",
   350 => x"ff497387",
   351 => x"7087cbdb",
   352 => x"c2c10298",
   353 => x"fd4cc187",
   354 => x"497587fd",
   355 => x"7087e3ca",
   356 => x"87c60298",
   357 => x"48e4f7c2",
   358 => x"f7c250c1",
   359 => x"05bf97e4",
   360 => x"c287e4c0",
   361 => x"49bfedf7",
   362 => x"059966d0",
   363 => x"c287d6ff",
   364 => x"49bfe5f7",
   365 => x"059966d4",
   366 => x"7387caff",
   367 => x"c9daff49",
   368 => x"05987087",
   369 => x"7487fefe",
   370 => x"87d7fb48",
   371 => x"5c5b5e0e",
   372 => x"86f40e5d",
   373 => x"ec4c4dc0",
   374 => x"a6c47ebf",
   375 => x"f1f7c248",
   376 => x"1ec178bf",
   377 => x"49c71ec0",
   378 => x"c887cafd",
   379 => x"02987086",
   380 => x"49ff87ce",
   381 => x"c187c7fb",
   382 => x"d9ff49da",
   383 => x"4dc187cc",
   384 => x"97e4f7c2",
   385 => x"87c302bf",
   386 => x"c287c0c9",
   387 => x"4bbfe9f7",
   388 => x"bfdee0c2",
   389 => x"87ebc005",
   390 => x"ff49fdc3",
   391 => x"c387ebd8",
   392 => x"d8ff49fa",
   393 => x"497387e4",
   394 => x"7199ffc3",
   395 => x"fb49c01e",
   396 => x"497387c6",
   397 => x"7129b7c8",
   398 => x"fa49c11e",
   399 => x"86c887fa",
   400 => x"c287c1c6",
   401 => x"4bbfedf7",
   402 => x"87dd029b",
   403 => x"bfdae0c2",
   404 => x"87dec749",
   405 => x"c4059870",
   406 => x"d24bc087",
   407 => x"49e0c287",
   408 => x"c287c3c7",
   409 => x"c658dee0",
   410 => x"dae0c287",
   411 => x"7378c048",
   412 => x"0599c249",
   413 => x"ebc387ce",
   414 => x"cdd7ff49",
   415 => x"c2497087",
   416 => x"87c20299",
   417 => x"49734cfb",
   418 => x"ce0599c1",
   419 => x"49f4c387",
   420 => x"87f6d6ff",
   421 => x"99c24970",
   422 => x"fa87c202",
   423 => x"c849734c",
   424 => x"87ce0599",
   425 => x"ff49f5c3",
   426 => x"7087dfd6",
   427 => x"0299c249",
   428 => x"f7c287d5",
   429 => x"ca02bff5",
   430 => x"88c14887",
   431 => x"58f9f7c2",
   432 => x"ff87c2c0",
   433 => x"734dc14c",
   434 => x"0599c449",
   435 => x"f2c387ce",
   436 => x"f5d5ff49",
   437 => x"c2497087",
   438 => x"87dc0299",
   439 => x"bff5f7c2",
   440 => x"b7c7487e",
   441 => x"cbc003a8",
   442 => x"c1486e87",
   443 => x"f9f7c280",
   444 => x"87c2c058",
   445 => x"4dc14cfe",
   446 => x"ff49fdc3",
   447 => x"7087cbd5",
   448 => x"0299c249",
   449 => x"c287d5c0",
   450 => x"02bff5f7",
   451 => x"c287c9c0",
   452 => x"c048f5f7",
   453 => x"87c2c078",
   454 => x"4dc14cfd",
   455 => x"ff49fac3",
   456 => x"7087e7d4",
   457 => x"0299c249",
   458 => x"c287d9c0",
   459 => x"48bff5f7",
   460 => x"03a8b7c7",
   461 => x"c287c9c0",
   462 => x"c748f5f7",
   463 => x"87c2c078",
   464 => x"4dc14cfc",
   465 => x"03acb7c0",
   466 => x"c487d1c0",
   467 => x"d8c14a66",
   468 => x"c0026a82",
   469 => x"4b6a87c6",
   470 => x"0f734974",
   471 => x"f0c31ec0",
   472 => x"49dac11e",
   473 => x"c887cef7",
   474 => x"02987086",
   475 => x"c887e2c0",
   476 => x"f7c248a6",
   477 => x"c878bff5",
   478 => x"91cb4966",
   479 => x"714866c4",
   480 => x"6e7e7080",
   481 => x"c8c002bf",
   482 => x"4bbf6e87",
   483 => x"734966c8",
   484 => x"029d750f",
   485 => x"c287c8c0",
   486 => x"49bff5f7",
   487 => x"c287faf2",
   488 => x"02bfe2e0",
   489 => x"4987ddc0",
   490 => x"7087c7c2",
   491 => x"d3c00298",
   492 => x"f5f7c287",
   493 => x"e0f249bf",
   494 => x"f449c087",
   495 => x"e0c287c0",
   496 => x"78c048e2",
   497 => x"daf38ef4",
   498 => x"5b5e0e87",
   499 => x"1e0e5d5c",
   500 => x"f7c24c71",
   501 => x"c149bff1",
   502 => x"c14da1cd",
   503 => x"7e6981d1",
   504 => x"cf029c74",
   505 => x"4ba5c487",
   506 => x"f7c27b74",
   507 => x"f249bff1",
   508 => x"7b6e87f9",
   509 => x"c4059c74",
   510 => x"c24bc087",
   511 => x"734bc187",
   512 => x"87faf249",
   513 => x"c70266d4",
   514 => x"87da4987",
   515 => x"87c24a70",
   516 => x"e0c24ac0",
   517 => x"f2265ae6",
   518 => x"000087c9",
   519 => x"00000000",
   520 => x"00000000",
   521 => x"711e0000",
   522 => x"bfc8ff4a",
   523 => x"48a17249",
   524 => x"ff1e4f26",
   525 => x"fe89bfc8",
   526 => x"c0c0c0c0",
   527 => x"c401a9c0",
   528 => x"c24ac087",
   529 => x"724ac187",
   530 => x"1e4f2648",
   531 => x"bfd9e2c2",
   532 => x"c2b9c149",
   533 => x"ff59dde2",
   534 => x"ffc348d4",
   535 => x"48d0ff78",
   536 => x"ff78e1c0",
   537 => x"78c148d4",
   538 => x"787131c4",
   539 => x"c048d0ff",
   540 => x"4f2678e0",
   541 => x"cde2c21e",
   542 => x"d8f2c21e",
   543 => x"c4fcfd49",
   544 => x"7086c487",
   545 => x"87c30298",
   546 => x"2687c0ff",
   547 => x"4b35314f",
   548 => x"20205a48",
   549 => x"47464320",
   550 => x"00000000",
   551 => x"5b5e0e00",
   552 => x"c20e5d5c",
   553 => x"4abfe5f7",
   554 => x"bfc6e4c2",
   555 => x"bc724c49",
   556 => x"c6ff4d71",
   557 => x"4bc087eb",
   558 => x"99d04974",
   559 => x"87e7c002",
   560 => x"c848d0ff",
   561 => x"d4ff78e1",
   562 => x"7578c548",
   563 => x"0299d049",
   564 => x"f0c387c3",
   565 => x"f4e4c278",
   566 => x"11817349",
   567 => x"08d4ff48",
   568 => x"48d0ff78",
   569 => x"c178e0c0",
   570 => x"c8832d2c",
   571 => x"c7ff04ab",
   572 => x"e4c5ff87",
   573 => x"c6e4c287",
   574 => x"e5f7c248",
   575 => x"4d2678bf",
   576 => x"4b264c26",
   577 => x"00004f26",
   578 => x"c11e0000",
   579 => x"de48cce7",
   580 => x"dde4c250",
   581 => x"f1d9fe49",
   582 => x"2648c087",
   583 => x"4f544a4f",
   584 => x"55525455",
   585 => x"4352414e",
   586 => x"dff21e00",
   587 => x"87edfd87",
   588 => x"4f2687f8",
   589 => x"25261e16",
   590 => x"3e3d362e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
