
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"ec",x"00",x"00",x"1f"),
     1 => (x"f1",x"00",x"00",x"1f"),
     2 => (x"1e",x"00",x"00",x"1f"),
     3 => (x"c8",x"48",x"d0",x"ff"),
     4 => (x"48",x"71",x"78",x"c9"),
     5 => (x"78",x"08",x"d4",x"ff"),
     6 => (x"71",x"1e",x"4f",x"26"),
     7 => (x"87",x"eb",x"49",x"4a"),
     8 => (x"c8",x"48",x"d0",x"ff"),
     9 => (x"1e",x"4f",x"26",x"78"),
    10 => (x"4b",x"71",x"1e",x"73"),
    11 => (x"bf",x"e4",x"f7",x"c2"),
    12 => (x"c2",x"87",x"c3",x"02"),
    13 => (x"d0",x"ff",x"87",x"eb"),
    14 => (x"78",x"c9",x"c8",x"48"),
    15 => (x"e0",x"c0",x"49",x"73"),
    16 => (x"48",x"d4",x"ff",x"b1"),
    17 => (x"f7",x"c2",x"78",x"71"),
    18 => (x"78",x"c0",x"48",x"d8"),
    19 => (x"c5",x"02",x"66",x"c8"),
    20 => (x"49",x"ff",x"c3",x"87"),
    21 => (x"49",x"c0",x"87",x"c2"),
    22 => (x"59",x"e0",x"f7",x"c2"),
    23 => (x"c6",x"02",x"66",x"cc"),
    24 => (x"d5",x"d5",x"c5",x"87"),
    25 => (x"cf",x"87",x"c4",x"4a"),
    26 => (x"c2",x"4a",x"ff",x"ff"),
    27 => (x"c2",x"5a",x"e4",x"f7"),
    28 => (x"c1",x"48",x"e4",x"f7"),
    29 => (x"26",x"87",x"c4",x"78"),
    30 => (x"26",x"4c",x"26",x"4d"),
    31 => (x"0e",x"4f",x"26",x"4b"),
    32 => (x"5d",x"5c",x"5b",x"5e"),
    33 => (x"c2",x"4a",x"71",x"0e"),
    34 => (x"4c",x"bf",x"e0",x"f7"),
    35 => (x"cb",x"02",x"9a",x"72"),
    36 => (x"91",x"c8",x"49",x"87"),
    37 => (x"4b",x"dd",x"c0",x"c2"),
    38 => (x"87",x"c4",x"83",x"71"),
    39 => (x"4b",x"dd",x"c4",x"c2"),
    40 => (x"49",x"13",x"4d",x"c0"),
    41 => (x"f7",x"c2",x"99",x"74"),
    42 => (x"ff",x"b9",x"bf",x"dc"),
    43 => (x"78",x"71",x"48",x"d4"),
    44 => (x"85",x"2c",x"b7",x"c1"),
    45 => (x"04",x"ad",x"b7",x"c8"),
    46 => (x"f7",x"c2",x"87",x"e8"),
    47 => (x"c8",x"48",x"bf",x"d8"),
    48 => (x"dc",x"f7",x"c2",x"80"),
    49 => (x"87",x"ef",x"fe",x"58"),
    50 => (x"71",x"1e",x"73",x"1e"),
    51 => (x"9a",x"4a",x"13",x"4b"),
    52 => (x"72",x"87",x"cb",x"02"),
    53 => (x"87",x"e7",x"fe",x"49"),
    54 => (x"05",x"9a",x"4a",x"13"),
    55 => (x"da",x"fe",x"87",x"f5"),
    56 => (x"f7",x"c2",x"1e",x"87"),
    57 => (x"c2",x"49",x"bf",x"d8"),
    58 => (x"c1",x"48",x"d8",x"f7"),
    59 => (x"c0",x"c4",x"78",x"a1"),
    60 => (x"db",x"03",x"a9",x"b7"),
    61 => (x"48",x"d4",x"ff",x"87"),
    62 => (x"bf",x"dc",x"f7",x"c2"),
    63 => (x"d8",x"f7",x"c2",x"78"),
    64 => (x"f7",x"c2",x"49",x"bf"),
    65 => (x"a1",x"c1",x"48",x"d8"),
    66 => (x"b7",x"c0",x"c4",x"78"),
    67 => (x"87",x"e5",x"04",x"a9"),
    68 => (x"c8",x"48",x"d0",x"ff"),
    69 => (x"e4",x"f7",x"c2",x"78"),
    70 => (x"26",x"78",x"c0",x"48"),
    71 => (x"00",x"00",x"00",x"4f"),
    72 => (x"00",x"00",x"00",x"00"),
    73 => (x"00",x"00",x"00",x"00"),
    74 => (x"00",x"00",x"5f",x"5f"),
    75 => (x"03",x"03",x"00",x"00"),
    76 => (x"00",x"03",x"03",x"00"),
    77 => (x"7f",x"7f",x"14",x"00"),
    78 => (x"14",x"7f",x"7f",x"14"),
    79 => (x"2e",x"24",x"00",x"00"),
    80 => (x"12",x"3a",x"6b",x"6b"),
    81 => (x"36",x"6a",x"4c",x"00"),
    82 => (x"32",x"56",x"6c",x"18"),
    83 => (x"4f",x"7e",x"30",x"00"),
    84 => (x"68",x"3a",x"77",x"59"),
    85 => (x"04",x"00",x"00",x"40"),
    86 => (x"00",x"00",x"03",x"07"),
    87 => (x"1c",x"00",x"00",x"00"),
    88 => (x"00",x"41",x"63",x"3e"),
    89 => (x"41",x"00",x"00",x"00"),
    90 => (x"00",x"1c",x"3e",x"63"),
    91 => (x"3e",x"2a",x"08",x"00"),
    92 => (x"2a",x"3e",x"1c",x"1c"),
    93 => (x"08",x"08",x"00",x"08"),
    94 => (x"08",x"08",x"3e",x"3e"),
    95 => (x"80",x"00",x"00",x"00"),
    96 => (x"00",x"00",x"60",x"e0"),
    97 => (x"08",x"08",x"00",x"00"),
    98 => (x"08",x"08",x"08",x"08"),
    99 => (x"00",x"00",x"00",x"00"),
   100 => (x"00",x"00",x"60",x"60"),
   101 => (x"30",x"60",x"40",x"00"),
   102 => (x"03",x"06",x"0c",x"18"),
   103 => (x"7f",x"3e",x"00",x"01"),
   104 => (x"3e",x"7f",x"4d",x"59"),
   105 => (x"06",x"04",x"00",x"00"),
   106 => (x"00",x"00",x"7f",x"7f"),
   107 => (x"63",x"42",x"00",x"00"),
   108 => (x"46",x"4f",x"59",x"71"),
   109 => (x"63",x"22",x"00",x"00"),
   110 => (x"36",x"7f",x"49",x"49"),
   111 => (x"16",x"1c",x"18",x"00"),
   112 => (x"10",x"7f",x"7f",x"13"),
   113 => (x"67",x"27",x"00",x"00"),
   114 => (x"39",x"7d",x"45",x"45"),
   115 => (x"7e",x"3c",x"00",x"00"),
   116 => (x"30",x"79",x"49",x"4b"),
   117 => (x"01",x"01",x"00",x"00"),
   118 => (x"07",x"0f",x"79",x"71"),
   119 => (x"7f",x"36",x"00",x"00"),
   120 => (x"36",x"7f",x"49",x"49"),
   121 => (x"4f",x"06",x"00",x"00"),
   122 => (x"1e",x"3f",x"69",x"49"),
   123 => (x"00",x"00",x"00",x"00"),
   124 => (x"00",x"00",x"66",x"66"),
   125 => (x"80",x"00",x"00",x"00"),
   126 => (x"00",x"00",x"66",x"e6"),
   127 => (x"08",x"08",x"00",x"00"),
   128 => (x"22",x"22",x"14",x"14"),
   129 => (x"14",x"14",x"00",x"00"),
   130 => (x"14",x"14",x"14",x"14"),
   131 => (x"22",x"22",x"00",x"00"),
   132 => (x"08",x"08",x"14",x"14"),
   133 => (x"03",x"02",x"00",x"00"),
   134 => (x"06",x"0f",x"59",x"51"),
   135 => (x"41",x"7f",x"3e",x"00"),
   136 => (x"1e",x"1f",x"55",x"5d"),
   137 => (x"7f",x"7e",x"00",x"00"),
   138 => (x"7e",x"7f",x"09",x"09"),
   139 => (x"7f",x"7f",x"00",x"00"),
   140 => (x"36",x"7f",x"49",x"49"),
   141 => (x"3e",x"1c",x"00",x"00"),
   142 => (x"41",x"41",x"41",x"63"),
   143 => (x"7f",x"7f",x"00",x"00"),
   144 => (x"1c",x"3e",x"63",x"41"),
   145 => (x"7f",x"7f",x"00",x"00"),
   146 => (x"41",x"41",x"49",x"49"),
   147 => (x"7f",x"7f",x"00",x"00"),
   148 => (x"01",x"01",x"09",x"09"),
   149 => (x"7f",x"3e",x"00",x"00"),
   150 => (x"7a",x"7b",x"49",x"41"),
   151 => (x"7f",x"7f",x"00",x"00"),
   152 => (x"7f",x"7f",x"08",x"08"),
   153 => (x"41",x"00",x"00",x"00"),
   154 => (x"00",x"41",x"7f",x"7f"),
   155 => (x"60",x"20",x"00",x"00"),
   156 => (x"3f",x"7f",x"40",x"40"),
   157 => (x"08",x"7f",x"7f",x"00"),
   158 => (x"41",x"63",x"36",x"1c"),
   159 => (x"7f",x"7f",x"00",x"00"),
   160 => (x"40",x"40",x"40",x"40"),
   161 => (x"06",x"7f",x"7f",x"00"),
   162 => (x"7f",x"7f",x"06",x"0c"),
   163 => (x"06",x"7f",x"7f",x"00"),
   164 => (x"7f",x"7f",x"18",x"0c"),
   165 => (x"7f",x"3e",x"00",x"00"),
   166 => (x"3e",x"7f",x"41",x"41"),
   167 => (x"7f",x"7f",x"00",x"00"),
   168 => (x"06",x"0f",x"09",x"09"),
   169 => (x"41",x"7f",x"3e",x"00"),
   170 => (x"40",x"7e",x"7f",x"61"),
   171 => (x"7f",x"7f",x"00",x"00"),
   172 => (x"66",x"7f",x"19",x"09"),
   173 => (x"6f",x"26",x"00",x"00"),
   174 => (x"32",x"7b",x"59",x"4d"),
   175 => (x"01",x"01",x"00",x"00"),
   176 => (x"01",x"01",x"7f",x"7f"),
   177 => (x"7f",x"3f",x"00",x"00"),
   178 => (x"3f",x"7f",x"40",x"40"),
   179 => (x"3f",x"0f",x"00",x"00"),
   180 => (x"0f",x"3f",x"70",x"70"),
   181 => (x"30",x"7f",x"7f",x"00"),
   182 => (x"7f",x"7f",x"30",x"18"),
   183 => (x"36",x"63",x"41",x"00"),
   184 => (x"63",x"36",x"1c",x"1c"),
   185 => (x"06",x"03",x"01",x"41"),
   186 => (x"03",x"06",x"7c",x"7c"),
   187 => (x"59",x"71",x"61",x"01"),
   188 => (x"41",x"43",x"47",x"4d"),
   189 => (x"7f",x"00",x"00",x"00"),
   190 => (x"00",x"41",x"41",x"7f"),
   191 => (x"06",x"03",x"01",x"00"),
   192 => (x"60",x"30",x"18",x"0c"),
   193 => (x"41",x"00",x"00",x"40"),
   194 => (x"00",x"7f",x"7f",x"41"),
   195 => (x"06",x"0c",x"08",x"00"),
   196 => (x"08",x"0c",x"06",x"03"),
   197 => (x"80",x"80",x"80",x"00"),
   198 => (x"80",x"80",x"80",x"80"),
   199 => (x"00",x"00",x"00",x"00"),
   200 => (x"00",x"04",x"07",x"03"),
   201 => (x"74",x"20",x"00",x"00"),
   202 => (x"78",x"7c",x"54",x"54"),
   203 => (x"7f",x"7f",x"00",x"00"),
   204 => (x"38",x"7c",x"44",x"44"),
   205 => (x"7c",x"38",x"00",x"00"),
   206 => (x"00",x"44",x"44",x"44"),
   207 => (x"7c",x"38",x"00",x"00"),
   208 => (x"7f",x"7f",x"44",x"44"),
   209 => (x"7c",x"38",x"00",x"00"),
   210 => (x"18",x"5c",x"54",x"54"),
   211 => (x"7e",x"04",x"00",x"00"),
   212 => (x"00",x"05",x"05",x"7f"),
   213 => (x"bc",x"18",x"00",x"00"),
   214 => (x"7c",x"fc",x"a4",x"a4"),
   215 => (x"7f",x"7f",x"00",x"00"),
   216 => (x"78",x"7c",x"04",x"04"),
   217 => (x"00",x"00",x"00",x"00"),
   218 => (x"00",x"40",x"7d",x"3d"),
   219 => (x"80",x"80",x"00",x"00"),
   220 => (x"00",x"7d",x"fd",x"80"),
   221 => (x"7f",x"7f",x"00",x"00"),
   222 => (x"44",x"6c",x"38",x"10"),
   223 => (x"00",x"00",x"00",x"00"),
   224 => (x"00",x"40",x"7f",x"3f"),
   225 => (x"0c",x"7c",x"7c",x"00"),
   226 => (x"78",x"7c",x"0c",x"18"),
   227 => (x"7c",x"7c",x"00",x"00"),
   228 => (x"78",x"7c",x"04",x"04"),
   229 => (x"7c",x"38",x"00",x"00"),
   230 => (x"38",x"7c",x"44",x"44"),
   231 => (x"fc",x"fc",x"00",x"00"),
   232 => (x"18",x"3c",x"24",x"24"),
   233 => (x"3c",x"18",x"00",x"00"),
   234 => (x"fc",x"fc",x"24",x"24"),
   235 => (x"7c",x"7c",x"00",x"00"),
   236 => (x"08",x"0c",x"04",x"04"),
   237 => (x"5c",x"48",x"00",x"00"),
   238 => (x"20",x"74",x"54",x"54"),
   239 => (x"3f",x"04",x"00",x"00"),
   240 => (x"00",x"44",x"44",x"7f"),
   241 => (x"7c",x"3c",x"00",x"00"),
   242 => (x"7c",x"7c",x"40",x"40"),
   243 => (x"3c",x"1c",x"00",x"00"),
   244 => (x"1c",x"3c",x"60",x"60"),
   245 => (x"60",x"7c",x"3c",x"00"),
   246 => (x"3c",x"7c",x"60",x"30"),
   247 => (x"38",x"6c",x"44",x"00"),
   248 => (x"44",x"6c",x"38",x"10"),
   249 => (x"bc",x"1c",x"00",x"00"),
   250 => (x"1c",x"3c",x"60",x"e0"),
   251 => (x"64",x"44",x"00",x"00"),
   252 => (x"44",x"4c",x"5c",x"74"),
   253 => (x"08",x"08",x"00",x"00"),
   254 => (x"41",x"41",x"77",x"3e"),
   255 => (x"00",x"00",x"00",x"00"),
   256 => (x"00",x"00",x"7f",x"7f"),
   257 => (x"41",x"41",x"00",x"00"),
   258 => (x"08",x"08",x"3e",x"77"),
   259 => (x"01",x"01",x"02",x"00"),
   260 => (x"01",x"02",x"02",x"03"),
   261 => (x"7f",x"7f",x"7f",x"00"),
   262 => (x"7f",x"7f",x"7f",x"7f"),
   263 => (x"1c",x"08",x"08",x"00"),
   264 => (x"7f",x"3e",x"3e",x"1c"),
   265 => (x"3e",x"7f",x"7f",x"7f"),
   266 => (x"08",x"1c",x"1c",x"3e"),
   267 => (x"18",x"10",x"00",x"08"),
   268 => (x"10",x"18",x"7c",x"7c"),
   269 => (x"30",x"10",x"00",x"00"),
   270 => (x"10",x"30",x"7c",x"7c"),
   271 => (x"60",x"30",x"10",x"00"),
   272 => (x"06",x"1e",x"78",x"60"),
   273 => (x"3c",x"66",x"42",x"00"),
   274 => (x"42",x"66",x"3c",x"18"),
   275 => (x"6a",x"38",x"78",x"00"),
   276 => (x"38",x"6c",x"c6",x"c2"),
   277 => (x"00",x"00",x"60",x"00"),
   278 => (x"60",x"00",x"00",x"60"),
   279 => (x"5b",x"5e",x"0e",x"00"),
   280 => (x"1e",x"0e",x"5d",x"5c"),
   281 => (x"f7",x"c2",x"4c",x"71"),
   282 => (x"c0",x"4d",x"bf",x"f5"),
   283 => (x"74",x"1e",x"c0",x"4b"),
   284 => (x"87",x"c7",x"02",x"ab"),
   285 => (x"c0",x"48",x"a6",x"c4"),
   286 => (x"c4",x"87",x"c5",x"78"),
   287 => (x"78",x"c1",x"48",x"a6"),
   288 => (x"73",x"1e",x"66",x"c4"),
   289 => (x"87",x"df",x"ee",x"49"),
   290 => (x"e0",x"c0",x"86",x"c8"),
   291 => (x"87",x"ef",x"ef",x"49"),
   292 => (x"6a",x"4a",x"a5",x"c4"),
   293 => (x"87",x"f0",x"f0",x"49"),
   294 => (x"cb",x"87",x"c6",x"f1"),
   295 => (x"c8",x"83",x"c1",x"85"),
   296 => (x"ff",x"04",x"ab",x"b7"),
   297 => (x"26",x"26",x"87",x"c7"),
   298 => (x"26",x"4c",x"26",x"4d"),
   299 => (x"1e",x"4f",x"26",x"4b"),
   300 => (x"f7",x"c2",x"4a",x"71"),
   301 => (x"f7",x"c2",x"5a",x"f9"),
   302 => (x"78",x"c7",x"48",x"f9"),
   303 => (x"87",x"dd",x"fe",x"49"),
   304 => (x"73",x"1e",x"4f",x"26"),
   305 => (x"c0",x"4a",x"71",x"1e"),
   306 => (x"d3",x"03",x"aa",x"b7"),
   307 => (x"e2",x"e0",x"c2",x"87"),
   308 => (x"87",x"c4",x"05",x"bf"),
   309 => (x"87",x"c2",x"4b",x"c1"),
   310 => (x"e0",x"c2",x"4b",x"c0"),
   311 => (x"87",x"c4",x"5b",x"e6"),
   312 => (x"5a",x"e6",x"e0",x"c2"),
   313 => (x"bf",x"e2",x"e0",x"c2"),
   314 => (x"c1",x"9a",x"c1",x"4a"),
   315 => (x"ec",x"49",x"a2",x"c0"),
   316 => (x"48",x"fc",x"87",x"e8"),
   317 => (x"bf",x"e2",x"e0",x"c2"),
   318 => (x"87",x"ef",x"fe",x"78"),
   319 => (x"c4",x"4a",x"71",x"1e"),
   320 => (x"49",x"72",x"1e",x"66"),
   321 => (x"87",x"e9",x"df",x"ff"),
   322 => (x"1e",x"4f",x"26",x"26"),
   323 => (x"bf",x"e2",x"e0",x"c2"),
   324 => (x"d9",x"dc",x"ff",x"49"),
   325 => (x"ed",x"f7",x"c2",x"87"),
   326 => (x"78",x"bf",x"e8",x"48"),
   327 => (x"48",x"e9",x"f7",x"c2"),
   328 => (x"c2",x"78",x"bf",x"ec"),
   329 => (x"4a",x"bf",x"ed",x"f7"),
   330 => (x"99",x"ff",x"c3",x"49"),
   331 => (x"72",x"2a",x"b7",x"c8"),
   332 => (x"c2",x"b0",x"71",x"48"),
   333 => (x"26",x"58",x"f5",x"f7"),
   334 => (x"5b",x"5e",x"0e",x"4f"),
   335 => (x"71",x"0e",x"5d",x"5c"),
   336 => (x"87",x"c7",x"ff",x"4b"),
   337 => (x"48",x"e8",x"f7",x"c2"),
   338 => (x"49",x"73",x"50",x"c0"),
   339 => (x"87",x"fe",x"db",x"ff"),
   340 => (x"c2",x"4c",x"49",x"70"),
   341 => (x"49",x"ee",x"cb",x"9c"),
   342 => (x"70",x"87",x"cf",x"cb"),
   343 => (x"f7",x"c2",x"4d",x"49"),
   344 => (x"05",x"bf",x"97",x"e8"),
   345 => (x"d0",x"87",x"e4",x"c1"),
   346 => (x"f7",x"c2",x"49",x"66"),
   347 => (x"05",x"99",x"bf",x"f1"),
   348 => (x"66",x"d4",x"87",x"d7"),
   349 => (x"e9",x"f7",x"c2",x"49"),
   350 => (x"cc",x"05",x"99",x"bf"),
   351 => (x"ff",x"49",x"73",x"87"),
   352 => (x"70",x"87",x"cb",x"db"),
   353 => (x"c2",x"c1",x"02",x"98"),
   354 => (x"fd",x"4c",x"c1",x"87"),
   355 => (x"49",x"75",x"87",x"fd"),
   356 => (x"70",x"87",x"e3",x"ca"),
   357 => (x"87",x"c6",x"02",x"98"),
   358 => (x"48",x"e8",x"f7",x"c2"),
   359 => (x"f7",x"c2",x"50",x"c1"),
   360 => (x"05",x"bf",x"97",x"e8"),
   361 => (x"c2",x"87",x"e4",x"c0"),
   362 => (x"49",x"bf",x"f1",x"f7"),
   363 => (x"05",x"99",x"66",x"d0"),
   364 => (x"c2",x"87",x"d6",x"ff"),
   365 => (x"49",x"bf",x"e9",x"f7"),
   366 => (x"05",x"99",x"66",x"d4"),
   367 => (x"73",x"87",x"ca",x"ff"),
   368 => (x"c9",x"da",x"ff",x"49"),
   369 => (x"05",x"98",x"70",x"87"),
   370 => (x"74",x"87",x"fe",x"fe"),
   371 => (x"87",x"d7",x"fb",x"48"),
   372 => (x"5c",x"5b",x"5e",x"0e"),
   373 => (x"86",x"f4",x"0e",x"5d"),
   374 => (x"ec",x"4c",x"4d",x"c0"),
   375 => (x"a6",x"c4",x"7e",x"bf"),
   376 => (x"f5",x"f7",x"c2",x"48"),
   377 => (x"1e",x"c1",x"78",x"bf"),
   378 => (x"49",x"c7",x"1e",x"c0"),
   379 => (x"c8",x"87",x"ca",x"fd"),
   380 => (x"02",x"98",x"70",x"86"),
   381 => (x"49",x"ff",x"87",x"ce"),
   382 => (x"c1",x"87",x"c7",x"fb"),
   383 => (x"d9",x"ff",x"49",x"da"),
   384 => (x"4d",x"c1",x"87",x"cc"),
   385 => (x"97",x"e8",x"f7",x"c2"),
   386 => (x"87",x"c3",x"02",x"bf"),
   387 => (x"c2",x"87",x"c0",x"c9"),
   388 => (x"4b",x"bf",x"ed",x"f7"),
   389 => (x"bf",x"e2",x"e0",x"c2"),
   390 => (x"87",x"eb",x"c0",x"05"),
   391 => (x"ff",x"49",x"fd",x"c3"),
   392 => (x"c3",x"87",x"eb",x"d8"),
   393 => (x"d8",x"ff",x"49",x"fa"),
   394 => (x"49",x"73",x"87",x"e4"),
   395 => (x"71",x"99",x"ff",x"c3"),
   396 => (x"fb",x"49",x"c0",x"1e"),
   397 => (x"49",x"73",x"87",x"c6"),
   398 => (x"71",x"29",x"b7",x"c8"),
   399 => (x"fa",x"49",x"c1",x"1e"),
   400 => (x"86",x"c8",x"87",x"fa"),
   401 => (x"c2",x"87",x"c1",x"c6"),
   402 => (x"4b",x"bf",x"f1",x"f7"),
   403 => (x"87",x"dd",x"02",x"9b"),
   404 => (x"bf",x"de",x"e0",x"c2"),
   405 => (x"87",x"de",x"c7",x"49"),
   406 => (x"c4",x"05",x"98",x"70"),
   407 => (x"d2",x"4b",x"c0",x"87"),
   408 => (x"49",x"e0",x"c2",x"87"),
   409 => (x"c2",x"87",x"c3",x"c7"),
   410 => (x"c6",x"58",x"e2",x"e0"),
   411 => (x"de",x"e0",x"c2",x"87"),
   412 => (x"73",x"78",x"c0",x"48"),
   413 => (x"05",x"99",x"c2",x"49"),
   414 => (x"eb",x"c3",x"87",x"ce"),
   415 => (x"cd",x"d7",x"ff",x"49"),
   416 => (x"c2",x"49",x"70",x"87"),
   417 => (x"87",x"c2",x"02",x"99"),
   418 => (x"49",x"73",x"4c",x"fb"),
   419 => (x"ce",x"05",x"99",x"c1"),
   420 => (x"49",x"f4",x"c3",x"87"),
   421 => (x"87",x"f6",x"d6",x"ff"),
   422 => (x"99",x"c2",x"49",x"70"),
   423 => (x"fa",x"87",x"c2",x"02"),
   424 => (x"c8",x"49",x"73",x"4c"),
   425 => (x"87",x"ce",x"05",x"99"),
   426 => (x"ff",x"49",x"f5",x"c3"),
   427 => (x"70",x"87",x"df",x"d6"),
   428 => (x"02",x"99",x"c2",x"49"),
   429 => (x"f7",x"c2",x"87",x"d5"),
   430 => (x"ca",x"02",x"bf",x"f9"),
   431 => (x"88",x"c1",x"48",x"87"),
   432 => (x"58",x"fd",x"f7",x"c2"),
   433 => (x"ff",x"87",x"c2",x"c0"),
   434 => (x"73",x"4d",x"c1",x"4c"),
   435 => (x"05",x"99",x"c4",x"49"),
   436 => (x"f2",x"c3",x"87",x"ce"),
   437 => (x"f5",x"d5",x"ff",x"49"),
   438 => (x"c2",x"49",x"70",x"87"),
   439 => (x"87",x"dc",x"02",x"99"),
   440 => (x"bf",x"f9",x"f7",x"c2"),
   441 => (x"b7",x"c7",x"48",x"7e"),
   442 => (x"cb",x"c0",x"03",x"a8"),
   443 => (x"c1",x"48",x"6e",x"87"),
   444 => (x"fd",x"f7",x"c2",x"80"),
   445 => (x"87",x"c2",x"c0",x"58"),
   446 => (x"4d",x"c1",x"4c",x"fe"),
   447 => (x"ff",x"49",x"fd",x"c3"),
   448 => (x"70",x"87",x"cb",x"d5"),
   449 => (x"02",x"99",x"c2",x"49"),
   450 => (x"c2",x"87",x"d5",x"c0"),
   451 => (x"02",x"bf",x"f9",x"f7"),
   452 => (x"c2",x"87",x"c9",x"c0"),
   453 => (x"c0",x"48",x"f9",x"f7"),
   454 => (x"87",x"c2",x"c0",x"78"),
   455 => (x"4d",x"c1",x"4c",x"fd"),
   456 => (x"ff",x"49",x"fa",x"c3"),
   457 => (x"70",x"87",x"e7",x"d4"),
   458 => (x"02",x"99",x"c2",x"49"),
   459 => (x"c2",x"87",x"d9",x"c0"),
   460 => (x"48",x"bf",x"f9",x"f7"),
   461 => (x"03",x"a8",x"b7",x"c7"),
   462 => (x"c2",x"87",x"c9",x"c0"),
   463 => (x"c7",x"48",x"f9",x"f7"),
   464 => (x"87",x"c2",x"c0",x"78"),
   465 => (x"4d",x"c1",x"4c",x"fc"),
   466 => (x"03",x"ac",x"b7",x"c0"),
   467 => (x"c4",x"87",x"d1",x"c0"),
   468 => (x"d8",x"c1",x"4a",x"66"),
   469 => (x"c0",x"02",x"6a",x"82"),
   470 => (x"4b",x"6a",x"87",x"c6"),
   471 => (x"0f",x"73",x"49",x"74"),
   472 => (x"f0",x"c3",x"1e",x"c0"),
   473 => (x"49",x"da",x"c1",x"1e"),
   474 => (x"c8",x"87",x"ce",x"f7"),
   475 => (x"02",x"98",x"70",x"86"),
   476 => (x"c8",x"87",x"e2",x"c0"),
   477 => (x"f7",x"c2",x"48",x"a6"),
   478 => (x"c8",x"78",x"bf",x"f9"),
   479 => (x"91",x"cb",x"49",x"66"),
   480 => (x"71",x"48",x"66",x"c4"),
   481 => (x"6e",x"7e",x"70",x"80"),
   482 => (x"c8",x"c0",x"02",x"bf"),
   483 => (x"4b",x"bf",x"6e",x"87"),
   484 => (x"73",x"49",x"66",x"c8"),
   485 => (x"02",x"9d",x"75",x"0f"),
   486 => (x"c2",x"87",x"c8",x"c0"),
   487 => (x"49",x"bf",x"f9",x"f7"),
   488 => (x"c2",x"87",x"fa",x"f2"),
   489 => (x"02",x"bf",x"e6",x"e0"),
   490 => (x"49",x"87",x"dd",x"c0"),
   491 => (x"70",x"87",x"c7",x"c2"),
   492 => (x"d3",x"c0",x"02",x"98"),
   493 => (x"f9",x"f7",x"c2",x"87"),
   494 => (x"e0",x"f2",x"49",x"bf"),
   495 => (x"f4",x"49",x"c0",x"87"),
   496 => (x"e0",x"c2",x"87",x"c0"),
   497 => (x"78",x"c0",x"48",x"e6"),
   498 => (x"da",x"f3",x"8e",x"f4"),
   499 => (x"5b",x"5e",x"0e",x"87"),
   500 => (x"1e",x"0e",x"5d",x"5c"),
   501 => (x"f7",x"c2",x"4c",x"71"),
   502 => (x"c1",x"49",x"bf",x"f5"),
   503 => (x"c1",x"4d",x"a1",x"cd"),
   504 => (x"7e",x"69",x"81",x"d1"),
   505 => (x"cf",x"02",x"9c",x"74"),
   506 => (x"4b",x"a5",x"c4",x"87"),
   507 => (x"f7",x"c2",x"7b",x"74"),
   508 => (x"f2",x"49",x"bf",x"f5"),
   509 => (x"7b",x"6e",x"87",x"f9"),
   510 => (x"c4",x"05",x"9c",x"74"),
   511 => (x"c2",x"4b",x"c0",x"87"),
   512 => (x"73",x"4b",x"c1",x"87"),
   513 => (x"87",x"fa",x"f2",x"49"),
   514 => (x"c7",x"02",x"66",x"d4"),
   515 => (x"87",x"da",x"49",x"87"),
   516 => (x"87",x"c2",x"4a",x"70"),
   517 => (x"e0",x"c2",x"4a",x"c0"),
   518 => (x"f2",x"26",x"5a",x"ea"),
   519 => (x"00",x"00",x"87",x"c9"),
   520 => (x"00",x"00",x"00",x"00"),
   521 => (x"00",x"00",x"00",x"00"),
   522 => (x"71",x"1e",x"00",x"00"),
   523 => (x"bf",x"c8",x"ff",x"4a"),
   524 => (x"48",x"a1",x"72",x"49"),
   525 => (x"ff",x"1e",x"4f",x"26"),
   526 => (x"fe",x"89",x"bf",x"c8"),
   527 => (x"c0",x"c0",x"c0",x"c0"),
   528 => (x"c4",x"01",x"a9",x"c0"),
   529 => (x"c2",x"4a",x"c0",x"87"),
   530 => (x"72",x"4a",x"c1",x"87"),
   531 => (x"1e",x"4f",x"26",x"48"),
   532 => (x"bf",x"dd",x"e2",x"c2"),
   533 => (x"c2",x"b9",x"c1",x"49"),
   534 => (x"ff",x"59",x"e1",x"e2"),
   535 => (x"ff",x"c3",x"48",x"d4"),
   536 => (x"48",x"d0",x"ff",x"78"),
   537 => (x"ff",x"78",x"e1",x"c0"),
   538 => (x"78",x"c1",x"48",x"d4"),
   539 => (x"78",x"71",x"31",x"c4"),
   540 => (x"c0",x"48",x"d0",x"ff"),
   541 => (x"4f",x"26",x"78",x"e0"),
   542 => (x"d1",x"e2",x"c2",x"1e"),
   543 => (x"dc",x"f2",x"c2",x"1e"),
   544 => (x"c0",x"fc",x"fd",x"49"),
   545 => (x"70",x"86",x"c4",x"87"),
   546 => (x"87",x"c3",x"02",x"98"),
   547 => (x"26",x"87",x"c0",x"ff"),
   548 => (x"4b",x"35",x"31",x"4f"),
   549 => (x"20",x"20",x"5a",x"48"),
   550 => (x"47",x"46",x"43",x"20"),
   551 => (x"00",x"00",x"00",x"00"),
   552 => (x"5b",x"5e",x"0e",x"00"),
   553 => (x"c2",x"0e",x"5d",x"5c"),
   554 => (x"4a",x"bf",x"e9",x"f7"),
   555 => (x"bf",x"ca",x"e4",x"c2"),
   556 => (x"bc",x"72",x"4c",x"49"),
   557 => (x"c6",x"ff",x"4d",x"71"),
   558 => (x"4b",x"c0",x"87",x"eb"),
   559 => (x"99",x"d0",x"49",x"74"),
   560 => (x"87",x"e7",x"c0",x"02"),
   561 => (x"c8",x"48",x"d0",x"ff"),
   562 => (x"d4",x"ff",x"78",x"e1"),
   563 => (x"75",x"78",x"c5",x"48"),
   564 => (x"02",x"99",x"d0",x"49"),
   565 => (x"f0",x"c3",x"87",x"c3"),
   566 => (x"f8",x"e4",x"c2",x"78"),
   567 => (x"11",x"81",x"73",x"49"),
   568 => (x"08",x"d4",x"ff",x"48"),
   569 => (x"48",x"d0",x"ff",x"78"),
   570 => (x"c1",x"78",x"e0",x"c0"),
   571 => (x"c8",x"83",x"2d",x"2c"),
   572 => (x"c7",x"ff",x"04",x"ab"),
   573 => (x"e4",x"c5",x"ff",x"87"),
   574 => (x"ca",x"e4",x"c2",x"87"),
   575 => (x"e9",x"f7",x"c2",x"48"),
   576 => (x"4d",x"26",x"78",x"bf"),
   577 => (x"4b",x"26",x"4c",x"26"),
   578 => (x"00",x"00",x"4f",x"26"),
   579 => (x"c1",x"1e",x"00",x"00"),
   580 => (x"de",x"48",x"d0",x"e7"),
   581 => (x"e1",x"e4",x"c2",x"50"),
   582 => (x"f1",x"d9",x"fe",x"49"),
   583 => (x"26",x"48",x"c0",x"87"),
   584 => (x"4f",x"54",x"4a",x"4f"),
   585 => (x"55",x"52",x"54",x"55"),
   586 => (x"43",x"52",x"41",x"4e"),
   587 => (x"df",x"f2",x"1e",x"00"),
   588 => (x"87",x"ed",x"fd",x"87"),
   589 => (x"4f",x"26",x"87",x"f8"),
   590 => (x"25",x"26",x"1e",x"16"),
   591 => (x"3e",x"3d",x"36",x"2e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

