library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"5ca6c887",
     1 => x"03acb7c0",
     2 => x"4887c4c0",
     3 => x"c487cac0",
     4 => x"c6f90266",
     5 => x"ffc34887",
     6 => x"f88ef499",
     7 => x"4f4387cf",
     8 => x"003d464e",
     9 => x"00444f4d",
    10 => x"454d414e",
    11 => x"46454400",
    12 => x"544c5541",
    13 => x"1e00303d",
    14 => x"24000020",
    15 => x"28000020",
    16 => x"2d000020",
    17 => x"1e000020",
    18 => x"c848d0ff",
    19 => x"487178c9",
    20 => x"7808d4ff",
    21 => x"711e4f26",
    22 => x"87eb494a",
    23 => x"c848d0ff",
    24 => x"1e4f2678",
    25 => x"4b711e73",
    26 => x"bfe0f8c2",
    27 => x"c287c302",
    28 => x"d0ff87eb",
    29 => x"78c9c848",
    30 => x"e0c04973",
    31 => x"48d4ffb1",
    32 => x"f8c27871",
    33 => x"78c048d4",
    34 => x"c50266c8",
    35 => x"49ffc387",
    36 => x"49c087c2",
    37 => x"59dcf8c2",
    38 => x"c60266cc",
    39 => x"d5d5c587",
    40 => x"cf87c44a",
    41 => x"c24affff",
    42 => x"c25ae0f8",
    43 => x"c148e0f8",
    44 => x"2687c478",
    45 => x"264c264d",
    46 => x"0e4f264b",
    47 => x"5d5c5b5e",
    48 => x"c24a710e",
    49 => x"4cbfdcf8",
    50 => x"cb029a72",
    51 => x"91c84987",
    52 => x"4bd9c1c2",
    53 => x"87c48371",
    54 => x"4bd9c5c2",
    55 => x"49134dc0",
    56 => x"f8c29974",
    57 => x"ffb9bfd8",
    58 => x"787148d4",
    59 => x"852cb7c1",
    60 => x"04adb7c8",
    61 => x"f8c287e8",
    62 => x"c848bfd4",
    63 => x"d8f8c280",
    64 => x"87effe58",
    65 => x"711e731e",
    66 => x"9a4a134b",
    67 => x"7287cb02",
    68 => x"87e7fe49",
    69 => x"059a4a13",
    70 => x"dafe87f5",
    71 => x"f8c21e87",
    72 => x"c249bfd4",
    73 => x"c148d4f8",
    74 => x"c0c478a1",
    75 => x"db03a9b7",
    76 => x"48d4ff87",
    77 => x"bfd8f8c2",
    78 => x"d4f8c278",
    79 => x"f8c249bf",
    80 => x"a1c148d4",
    81 => x"b7c0c478",
    82 => x"87e504a9",
    83 => x"c848d0ff",
    84 => x"e0f8c278",
    85 => x"2678c048",
    86 => x"0000004f",
    87 => x"00000000",
    88 => x"00000000",
    89 => x"00005f5f",
    90 => x"03030000",
    91 => x"00030300",
    92 => x"7f7f1400",
    93 => x"147f7f14",
    94 => x"2e240000",
    95 => x"123a6b6b",
    96 => x"366a4c00",
    97 => x"32566c18",
    98 => x"4f7e3000",
    99 => x"683a7759",
   100 => x"04000040",
   101 => x"00000307",
   102 => x"1c000000",
   103 => x"0041633e",
   104 => x"41000000",
   105 => x"001c3e63",
   106 => x"3e2a0800",
   107 => x"2a3e1c1c",
   108 => x"08080008",
   109 => x"08083e3e",
   110 => x"80000000",
   111 => x"000060e0",
   112 => x"08080000",
   113 => x"08080808",
   114 => x"00000000",
   115 => x"00006060",
   116 => x"30604000",
   117 => x"03060c18",
   118 => x"7f3e0001",
   119 => x"3e7f4d59",
   120 => x"06040000",
   121 => x"00007f7f",
   122 => x"63420000",
   123 => x"464f5971",
   124 => x"63220000",
   125 => x"367f4949",
   126 => x"161c1800",
   127 => x"107f7f13",
   128 => x"67270000",
   129 => x"397d4545",
   130 => x"7e3c0000",
   131 => x"3079494b",
   132 => x"01010000",
   133 => x"070f7971",
   134 => x"7f360000",
   135 => x"367f4949",
   136 => x"4f060000",
   137 => x"1e3f6949",
   138 => x"00000000",
   139 => x"00006666",
   140 => x"80000000",
   141 => x"000066e6",
   142 => x"08080000",
   143 => x"22221414",
   144 => x"14140000",
   145 => x"14141414",
   146 => x"22220000",
   147 => x"08081414",
   148 => x"03020000",
   149 => x"060f5951",
   150 => x"417f3e00",
   151 => x"1e1f555d",
   152 => x"7f7e0000",
   153 => x"7e7f0909",
   154 => x"7f7f0000",
   155 => x"367f4949",
   156 => x"3e1c0000",
   157 => x"41414163",
   158 => x"7f7f0000",
   159 => x"1c3e6341",
   160 => x"7f7f0000",
   161 => x"41414949",
   162 => x"7f7f0000",
   163 => x"01010909",
   164 => x"7f3e0000",
   165 => x"7a7b4941",
   166 => x"7f7f0000",
   167 => x"7f7f0808",
   168 => x"41000000",
   169 => x"00417f7f",
   170 => x"60200000",
   171 => x"3f7f4040",
   172 => x"087f7f00",
   173 => x"4163361c",
   174 => x"7f7f0000",
   175 => x"40404040",
   176 => x"067f7f00",
   177 => x"7f7f060c",
   178 => x"067f7f00",
   179 => x"7f7f180c",
   180 => x"7f3e0000",
   181 => x"3e7f4141",
   182 => x"7f7f0000",
   183 => x"060f0909",
   184 => x"417f3e00",
   185 => x"407e7f61",
   186 => x"7f7f0000",
   187 => x"667f1909",
   188 => x"6f260000",
   189 => x"327b594d",
   190 => x"01010000",
   191 => x"01017f7f",
   192 => x"7f3f0000",
   193 => x"3f7f4040",
   194 => x"3f0f0000",
   195 => x"0f3f7070",
   196 => x"307f7f00",
   197 => x"7f7f3018",
   198 => x"36634100",
   199 => x"63361c1c",
   200 => x"06030141",
   201 => x"03067c7c",
   202 => x"59716101",
   203 => x"4143474d",
   204 => x"7f000000",
   205 => x"0041417f",
   206 => x"06030100",
   207 => x"6030180c",
   208 => x"41000040",
   209 => x"007f7f41",
   210 => x"060c0800",
   211 => x"080c0603",
   212 => x"80808000",
   213 => x"80808080",
   214 => x"00000000",
   215 => x"00040703",
   216 => x"74200000",
   217 => x"787c5454",
   218 => x"7f7f0000",
   219 => x"387c4444",
   220 => x"7c380000",
   221 => x"00444444",
   222 => x"7c380000",
   223 => x"7f7f4444",
   224 => x"7c380000",
   225 => x"185c5454",
   226 => x"7e040000",
   227 => x"0005057f",
   228 => x"bc180000",
   229 => x"7cfca4a4",
   230 => x"7f7f0000",
   231 => x"787c0404",
   232 => x"00000000",
   233 => x"00407d3d",
   234 => x"80800000",
   235 => x"007dfd80",
   236 => x"7f7f0000",
   237 => x"446c3810",
   238 => x"00000000",
   239 => x"00407f3f",
   240 => x"0c7c7c00",
   241 => x"787c0c18",
   242 => x"7c7c0000",
   243 => x"787c0404",
   244 => x"7c380000",
   245 => x"387c4444",
   246 => x"fcfc0000",
   247 => x"183c2424",
   248 => x"3c180000",
   249 => x"fcfc2424",
   250 => x"7c7c0000",
   251 => x"080c0404",
   252 => x"5c480000",
   253 => x"20745454",
   254 => x"3f040000",
   255 => x"0044447f",
   256 => x"7c3c0000",
   257 => x"7c7c4040",
   258 => x"3c1c0000",
   259 => x"1c3c6060",
   260 => x"607c3c00",
   261 => x"3c7c6030",
   262 => x"386c4400",
   263 => x"446c3810",
   264 => x"bc1c0000",
   265 => x"1c3c60e0",
   266 => x"64440000",
   267 => x"444c5c74",
   268 => x"08080000",
   269 => x"4141773e",
   270 => x"00000000",
   271 => x"00007f7f",
   272 => x"41410000",
   273 => x"08083e77",
   274 => x"01010200",
   275 => x"01020203",
   276 => x"7f7f7f00",
   277 => x"7f7f7f7f",
   278 => x"1c080800",
   279 => x"7f3e3e1c",
   280 => x"3e7f7f7f",
   281 => x"081c1c3e",
   282 => x"18100008",
   283 => x"10187c7c",
   284 => x"30100000",
   285 => x"10307c7c",
   286 => x"60301000",
   287 => x"061e7860",
   288 => x"3c664200",
   289 => x"42663c18",
   290 => x"6a387800",
   291 => x"386cc6c2",
   292 => x"00006000",
   293 => x"60000060",
   294 => x"5b5e0e00",
   295 => x"1e0e5d5c",
   296 => x"f8c24c71",
   297 => x"c04dbff1",
   298 => x"741ec04b",
   299 => x"87c702ab",
   300 => x"c048a6c4",
   301 => x"c487c578",
   302 => x"78c148a6",
   303 => x"731e66c4",
   304 => x"87dfee49",
   305 => x"e0c086c8",
   306 => x"87efef49",
   307 => x"6a4aa5c4",
   308 => x"87f0f049",
   309 => x"cb87c6f1",
   310 => x"c883c185",
   311 => x"ff04abb7",
   312 => x"262687c7",
   313 => x"264c264d",
   314 => x"1e4f264b",
   315 => x"f8c24a71",
   316 => x"f8c25af5",
   317 => x"78c748f5",
   318 => x"87ddfe49",
   319 => x"731e4f26",
   320 => x"c04a711e",
   321 => x"d303aab7",
   322 => x"dee1c287",
   323 => x"87c405bf",
   324 => x"87c24bc1",
   325 => x"e1c24bc0",
   326 => x"87c45be2",
   327 => x"5ae2e1c2",
   328 => x"bfdee1c2",
   329 => x"c19ac14a",
   330 => x"ec49a2c0",
   331 => x"48fc87e8",
   332 => x"bfdee1c2",
   333 => x"87effe78",
   334 => x"c44a711e",
   335 => x"49721e66",
   336 => x"87d2dfff",
   337 => x"1e4f2626",
   338 => x"bfdee1c2",
   339 => x"e5dbff49",
   340 => x"e9f8c287",
   341 => x"78bfe848",
   342 => x"48e5f8c2",
   343 => x"c278bfec",
   344 => x"4abfe9f8",
   345 => x"99ffc349",
   346 => x"722ab7c8",
   347 => x"c2b07148",
   348 => x"2658f1f8",
   349 => x"5b5e0e4f",
   350 => x"710e5d5c",
   351 => x"87c7ff4b",
   352 => x"48e4f8c2",
   353 => x"497350c0",
   354 => x"87cadbff",
   355 => x"c24c4970",
   356 => x"49eecb9c",
   357 => x"7087cfcb",
   358 => x"f8c24d49",
   359 => x"05bf97e4",
   360 => x"d087e4c1",
   361 => x"f8c24966",
   362 => x"0599bfed",
   363 => x"66d487d7",
   364 => x"e5f8c249",
   365 => x"cc0599bf",
   366 => x"ff497387",
   367 => x"7087d7da",
   368 => x"c2c10298",
   369 => x"fd4cc187",
   370 => x"497587fd",
   371 => x"7087e3ca",
   372 => x"87c60298",
   373 => x"48e4f8c2",
   374 => x"f8c250c1",
   375 => x"05bf97e4",
   376 => x"c287e4c0",
   377 => x"49bfedf8",
   378 => x"059966d0",
   379 => x"c287d6ff",
   380 => x"49bfe5f8",
   381 => x"059966d4",
   382 => x"7387caff",
   383 => x"d5d9ff49",
   384 => x"05987087",
   385 => x"7487fefe",
   386 => x"87d7fb48",
   387 => x"5c5b5e0e",
   388 => x"86f40e5d",
   389 => x"ec4c4dc0",
   390 => x"a6c47ebf",
   391 => x"f1f8c248",
   392 => x"1ec178bf",
   393 => x"49c71ec0",
   394 => x"c887cafd",
   395 => x"02987086",
   396 => x"49ff87ce",
   397 => x"c187c7fb",
   398 => x"d8ff49da",
   399 => x"4dc187d8",
   400 => x"97e4f8c2",
   401 => x"87c302bf",
   402 => x"c287c0c9",
   403 => x"4bbfe9f8",
   404 => x"bfdee1c2",
   405 => x"87ebc005",
   406 => x"ff49fdc3",
   407 => x"c387f7d7",
   408 => x"d7ff49fa",
   409 => x"497387f0",
   410 => x"7199ffc3",
   411 => x"fb49c01e",
   412 => x"497387c6",
   413 => x"7129b7c8",
   414 => x"fa49c11e",
   415 => x"86c887fa",
   416 => x"c287c1c6",
   417 => x"4bbfedf8",
   418 => x"87dd029b",
   419 => x"bfdae1c2",
   420 => x"87dec749",
   421 => x"c4059870",
   422 => x"d24bc087",
   423 => x"49e0c287",
   424 => x"c287c3c7",
   425 => x"c658dee1",
   426 => x"dae1c287",
   427 => x"7378c048",
   428 => x"0599c249",
   429 => x"ebc387ce",
   430 => x"d9d6ff49",
   431 => x"c2497087",
   432 => x"87c20299",
   433 => x"49734cfb",
   434 => x"ce0599c1",
   435 => x"49f4c387",
   436 => x"87c2d6ff",
   437 => x"99c24970",
   438 => x"fa87c202",
   439 => x"c849734c",
   440 => x"87ce0599",
   441 => x"ff49f5c3",
   442 => x"7087ebd5",
   443 => x"0299c249",
   444 => x"f8c287d5",
   445 => x"ca02bff5",
   446 => x"88c14887",
   447 => x"58f9f8c2",
   448 => x"ff87c2c0",
   449 => x"734dc14c",
   450 => x"0599c449",
   451 => x"f2c387ce",
   452 => x"c1d5ff49",
   453 => x"c2497087",
   454 => x"87dc0299",
   455 => x"bff5f8c2",
   456 => x"b7c7487e",
   457 => x"cbc003a8",
   458 => x"c1486e87",
   459 => x"f9f8c280",
   460 => x"87c2c058",
   461 => x"4dc14cfe",
   462 => x"ff49fdc3",
   463 => x"7087d7d4",
   464 => x"0299c249",
   465 => x"c287d5c0",
   466 => x"02bff5f8",
   467 => x"c287c9c0",
   468 => x"c048f5f8",
   469 => x"87c2c078",
   470 => x"4dc14cfd",
   471 => x"ff49fac3",
   472 => x"7087f3d3",
   473 => x"0299c249",
   474 => x"c287d9c0",
   475 => x"48bff5f8",
   476 => x"03a8b7c7",
   477 => x"c287c9c0",
   478 => x"c748f5f8",
   479 => x"87c2c078",
   480 => x"4dc14cfc",
   481 => x"03acb7c0",
   482 => x"c487d1c0",
   483 => x"d8c14a66",
   484 => x"c0026a82",
   485 => x"4b6a87c6",
   486 => x"0f734974",
   487 => x"f0c31ec0",
   488 => x"49dac11e",
   489 => x"c887cef7",
   490 => x"02987086",
   491 => x"c887e2c0",
   492 => x"f8c248a6",
   493 => x"c878bff5",
   494 => x"91cb4966",
   495 => x"714866c4",
   496 => x"6e7e7080",
   497 => x"c8c002bf",
   498 => x"4bbf6e87",
   499 => x"734966c8",
   500 => x"029d750f",
   501 => x"c287c8c0",
   502 => x"49bff5f8",
   503 => x"c287faf2",
   504 => x"02bfe2e1",
   505 => x"4987ddc0",
   506 => x"7087c7c2",
   507 => x"d3c00298",
   508 => x"f5f8c287",
   509 => x"e0f249bf",
   510 => x"f449c087",
   511 => x"e1c287c0",
   512 => x"78c048e2",
   513 => x"daf38ef4",
   514 => x"5b5e0e87",
   515 => x"1e0e5d5c",
   516 => x"f8c24c71",
   517 => x"c149bff1",
   518 => x"c14da1cd",
   519 => x"7e6981d1",
   520 => x"cf029c74",
   521 => x"4ba5c487",
   522 => x"f8c27b74",
   523 => x"f249bff1",
   524 => x"7b6e87f9",
   525 => x"c4059c74",
   526 => x"c24bc087",
   527 => x"734bc187",
   528 => x"87faf249",
   529 => x"c70266d4",
   530 => x"87da4987",
   531 => x"87c24a70",
   532 => x"e1c24ac0",
   533 => x"f2265ae6",
   534 => x"000087c9",
   535 => x"00000000",
   536 => x"00000000",
   537 => x"711e0000",
   538 => x"bfc8ff4a",
   539 => x"48a17249",
   540 => x"ff1e4f26",
   541 => x"fe89bfc8",
   542 => x"c0c0c0c0",
   543 => x"c401a9c0",
   544 => x"c24ac087",
   545 => x"724ac187",
   546 => x"1e4f2648",
   547 => x"bfd9e3c2",
   548 => x"c2b9c149",
   549 => x"ff59dde3",
   550 => x"ffc348d4",
   551 => x"48d0ff78",
   552 => x"ff78e1c0",
   553 => x"78c148d4",
   554 => x"787131c4",
   555 => x"c048d0ff",
   556 => x"4f2678e0",
   557 => x"cde3c21e",
   558 => x"d8f3c21e",
   559 => x"d1fbfd49",
   560 => x"7086c487",
   561 => x"87c30298",
   562 => x"2687c0ff",
   563 => x"4b35314f",
   564 => x"20205a48",
   565 => x"47464320",
   566 => x"00000000",
   567 => x"5b5e0e00",
   568 => x"c20e5d5c",
   569 => x"4abfe5f8",
   570 => x"bfc6e5c2",
   571 => x"bc724c49",
   572 => x"c5ff4d71",
   573 => x"4bc087f7",
   574 => x"99d04974",
   575 => x"87e7c002",
   576 => x"c848d0ff",
   577 => x"d4ff78e1",
   578 => x"7578c548",
   579 => x"0299d049",
   580 => x"f0c387c3",
   581 => x"f4e5c278",
   582 => x"11817349",
   583 => x"08d4ff48",
   584 => x"48d0ff78",
   585 => x"c178e0c0",
   586 => x"c8832d2c",
   587 => x"c7ff04ab",
   588 => x"f0c4ff87",
   589 => x"c6e5c287",
   590 => x"e5f8c248",
   591 => x"4d2678bf",
   592 => x"4b264c26",
   593 => x"00004f26",
   594 => x"c11e0000",
   595 => x"de48d0e7",
   596 => x"dde5c250",
   597 => x"fad8fe49",
   598 => x"2648c087",
   599 => x"4f544a4f",
   600 => x"55525455",
   601 => x"4352414e",
   602 => x"dff21e00",
   603 => x"87edfd87",
   604 => x"4f2687f8",
   605 => x"25261e16",
   606 => x"3e3d362e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
