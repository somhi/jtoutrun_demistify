library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e4fac287",
    12 => x"86c0c54e",
    13 => x"49e4fac2",
    14 => x"48d8e7c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087f4e5",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"711e4f26",
    53 => x"4966c44a",
    54 => x"c888c148",
    55 => x"997158a6",
    56 => x"ff87d602",
    57 => x"ffc348d4",
    58 => x"c4526878",
    59 => x"c1484966",
    60 => x"58a6c888",
    61 => x"ea059971",
    62 => x"1e4f2687",
    63 => x"d4ff1e73",
    64 => x"7bffc34b",
    65 => x"ffc34a6b",
    66 => x"c8496b7b",
    67 => x"c3b17232",
    68 => x"4a6b7bff",
    69 => x"b27131c8",
    70 => x"6b7bffc3",
    71 => x"7232c849",
    72 => x"c44871b1",
    73 => x"264d2687",
    74 => x"264b264c",
    75 => x"5b5e0e4f",
    76 => x"710e5d5c",
    77 => x"4cd4ff4a",
    78 => x"ffc34972",
    79 => x"c27c7199",
    80 => x"05bfd8e7",
    81 => x"66d087c8",
    82 => x"d430c948",
    83 => x"66d058a6",
    84 => x"c329d849",
    85 => x"7c7199ff",
    86 => x"d04966d0",
    87 => x"99ffc329",
    88 => x"66d07c71",
    89 => x"c329c849",
    90 => x"7c7199ff",
    91 => x"c34966d0",
    92 => x"7c7199ff",
    93 => x"29d04972",
    94 => x"7199ffc3",
    95 => x"c94b6c7c",
    96 => x"c34dfff0",
    97 => x"d005abff",
    98 => x"7cffc387",
    99 => x"8dc14b6c",
   100 => x"c387c602",
   101 => x"f002abff",
   102 => x"fe487387",
   103 => x"c01e87c7",
   104 => x"48d4ff49",
   105 => x"c178ffc3",
   106 => x"b7c8c381",
   107 => x"87f104a9",
   108 => x"731e4f26",
   109 => x"c487e71e",
   110 => x"c04bdff8",
   111 => x"f0ffc01e",
   112 => x"fd49f7c1",
   113 => x"86c487e7",
   114 => x"c005a8c1",
   115 => x"d4ff87ea",
   116 => x"78ffc348",
   117 => x"c0c0c0c1",
   118 => x"c01ec0c0",
   119 => x"e9c1f0e1",
   120 => x"87c9fd49",
   121 => x"987086c4",
   122 => x"ff87ca05",
   123 => x"ffc348d4",
   124 => x"cb48c178",
   125 => x"87e6fe87",
   126 => x"fe058bc1",
   127 => x"48c087fd",
   128 => x"1e87e6fc",
   129 => x"d4ff1e73",
   130 => x"78ffc348",
   131 => x"1ec04bd3",
   132 => x"c1f0ffc0",
   133 => x"d4fc49c1",
   134 => x"7086c487",
   135 => x"87ca0598",
   136 => x"c348d4ff",
   137 => x"48c178ff",
   138 => x"f1fd87cb",
   139 => x"058bc187",
   140 => x"c087dbff",
   141 => x"87f1fb48",
   142 => x"5c5b5e0e",
   143 => x"4cd4ff0e",
   144 => x"c687dbfd",
   145 => x"e1c01eea",
   146 => x"49c8c1f0",
   147 => x"c487defb",
   148 => x"02a8c186",
   149 => x"eafe87c8",
   150 => x"c148c087",
   151 => x"dafa87e2",
   152 => x"cf497087",
   153 => x"c699ffff",
   154 => x"c802a9ea",
   155 => x"87d3fe87",
   156 => x"cbc148c0",
   157 => x"7cffc387",
   158 => x"fc4bf1c0",
   159 => x"987087f4",
   160 => x"87ebc002",
   161 => x"ffc01ec0",
   162 => x"49fac1f0",
   163 => x"c487defa",
   164 => x"05987086",
   165 => x"ffc387d9",
   166 => x"c3496c7c",
   167 => x"7c7c7cff",
   168 => x"99c0c17c",
   169 => x"c187c402",
   170 => x"c087d548",
   171 => x"c287d148",
   172 => x"87c405ab",
   173 => x"87c848c0",
   174 => x"fe058bc1",
   175 => x"48c087fd",
   176 => x"1e87e4f9",
   177 => x"e7c21e73",
   178 => x"78c148d8",
   179 => x"d0ff4bc7",
   180 => x"fb78c248",
   181 => x"d0ff87c8",
   182 => x"c078c348",
   183 => x"d0e5c01e",
   184 => x"f949c0c1",
   185 => x"86c487c7",
   186 => x"c105a8c1",
   187 => x"abc24b87",
   188 => x"c087c505",
   189 => x"87f9c048",
   190 => x"ff058bc1",
   191 => x"f7fc87d0",
   192 => x"dce7c287",
   193 => x"05987058",
   194 => x"1ec187cd",
   195 => x"c1f0ffc0",
   196 => x"d8f849d0",
   197 => x"ff86c487",
   198 => x"ffc348d4",
   199 => x"87fcc278",
   200 => x"58e0e7c2",
   201 => x"c248d0ff",
   202 => x"48d4ff78",
   203 => x"c178ffc3",
   204 => x"87f5f748",
   205 => x"5c5b5e0e",
   206 => x"4b710e5d",
   207 => x"eec54cc0",
   208 => x"ff4adfcd",
   209 => x"ffc348d4",
   210 => x"c3496878",
   211 => x"c005a9fe",
   212 => x"4d7087fd",
   213 => x"cc029b73",
   214 => x"1e66d087",
   215 => x"f1f54973",
   216 => x"d686c487",
   217 => x"48d0ff87",
   218 => x"c378d1c4",
   219 => x"66d07dff",
   220 => x"d488c148",
   221 => x"987058a6",
   222 => x"ff87f005",
   223 => x"ffc348d4",
   224 => x"9b737878",
   225 => x"ff87c505",
   226 => x"78d048d0",
   227 => x"c14c4ac1",
   228 => x"eefe058a",
   229 => x"f6487487",
   230 => x"731e87cb",
   231 => x"c04a711e",
   232 => x"48d4ff4b",
   233 => x"ff78ffc3",
   234 => x"c3c448d0",
   235 => x"48d4ff78",
   236 => x"7278ffc3",
   237 => x"f0ffc01e",
   238 => x"f549d1c1",
   239 => x"86c487ef",
   240 => x"d2059870",
   241 => x"1ec0c887",
   242 => x"fd4966cc",
   243 => x"86c487e6",
   244 => x"d0ff4b70",
   245 => x"7378c248",
   246 => x"87cdf548",
   247 => x"5c5b5e0e",
   248 => x"1ec00e5d",
   249 => x"c1f0ffc0",
   250 => x"c0f549c9",
   251 => x"c21ed287",
   252 => x"fc49e0e7",
   253 => x"86c887fe",
   254 => x"84c14cc0",
   255 => x"04acb7d2",
   256 => x"e7c287f8",
   257 => x"49bf97e0",
   258 => x"c199c0c3",
   259 => x"c005a9c0",
   260 => x"e7c287e7",
   261 => x"49bf97e7",
   262 => x"e7c231d0",
   263 => x"4abf97e8",
   264 => x"b17232c8",
   265 => x"97e9e7c2",
   266 => x"71b14abf",
   267 => x"ffffcf4c",
   268 => x"84c19cff",
   269 => x"e7c134ca",
   270 => x"e9e7c287",
   271 => x"c149bf97",
   272 => x"c299c631",
   273 => x"bf97eae7",
   274 => x"2ab7c74a",
   275 => x"e7c2b172",
   276 => x"4abf97e5",
   277 => x"c29dcf4d",
   278 => x"bf97e6e7",
   279 => x"ca9ac34a",
   280 => x"e7e7c232",
   281 => x"c24bbf97",
   282 => x"c2b27333",
   283 => x"bf97e8e7",
   284 => x"9bc0c34b",
   285 => x"732bb7c6",
   286 => x"c181c2b2",
   287 => x"70307148",
   288 => x"7548c149",
   289 => x"724d7030",
   290 => x"7184c14c",
   291 => x"b7c0c894",
   292 => x"87cc06ad",
   293 => x"2db734c1",
   294 => x"adb7c0c8",
   295 => x"87f4ff01",
   296 => x"c0f24874",
   297 => x"5b5e0e87",
   298 => x"f80e5d5c",
   299 => x"c6f0c286",
   300 => x"c278c048",
   301 => x"c01efee7",
   302 => x"87defb49",
   303 => x"987086c4",
   304 => x"c087c505",
   305 => x"87cec948",
   306 => x"7ec14dc0",
   307 => x"bfe2f5c0",
   308 => x"f4e8c249",
   309 => x"4bc8714a",
   310 => x"7087cfee",
   311 => x"87c20598",
   312 => x"f5c07ec0",
   313 => x"c249bfde",
   314 => x"714ad0e9",
   315 => x"f9ed4bc8",
   316 => x"05987087",
   317 => x"7ec087c2",
   318 => x"fdc0026e",
   319 => x"c4efc287",
   320 => x"efc24dbf",
   321 => x"7ebf9ffc",
   322 => x"ead6c548",
   323 => x"87c705a8",
   324 => x"bfc4efc2",
   325 => x"6e87ce4d",
   326 => x"d5e9ca48",
   327 => x"87c502a8",
   328 => x"f1c748c0",
   329 => x"fee7c287",
   330 => x"f949751e",
   331 => x"86c487ec",
   332 => x"c5059870",
   333 => x"c748c087",
   334 => x"f5c087dc",
   335 => x"c249bfde",
   336 => x"714ad0e9",
   337 => x"e1ec4bc8",
   338 => x"05987087",
   339 => x"f0c287c8",
   340 => x"78c148c6",
   341 => x"f5c087da",
   342 => x"c249bfe2",
   343 => x"714af4e8",
   344 => x"c5ec4bc8",
   345 => x"02987087",
   346 => x"c087c5c0",
   347 => x"87e6c648",
   348 => x"97fcefc2",
   349 => x"d5c149bf",
   350 => x"cdc005a9",
   351 => x"fdefc287",
   352 => x"c249bf97",
   353 => x"c002a9ea",
   354 => x"48c087c5",
   355 => x"c287c7c6",
   356 => x"bf97fee7",
   357 => x"e9c3487e",
   358 => x"cec002a8",
   359 => x"c3486e87",
   360 => x"c002a8eb",
   361 => x"48c087c5",
   362 => x"c287ebc5",
   363 => x"bf97c9e8",
   364 => x"c0059949",
   365 => x"e8c287cc",
   366 => x"49bf97ca",
   367 => x"c002a9c2",
   368 => x"48c087c5",
   369 => x"c287cfc5",
   370 => x"bf97cbe8",
   371 => x"c2f0c248",
   372 => x"484c7058",
   373 => x"f0c288c1",
   374 => x"e8c258c6",
   375 => x"49bf97cc",
   376 => x"e8c28175",
   377 => x"4abf97cd",
   378 => x"a17232c8",
   379 => x"d3f4c27e",
   380 => x"c2786e48",
   381 => x"bf97cee8",
   382 => x"58a6c848",
   383 => x"bfc6f0c2",
   384 => x"87d4c202",
   385 => x"bfdef5c0",
   386 => x"d0e9c249",
   387 => x"4bc8714a",
   388 => x"7087d7e9",
   389 => x"c5c00298",
   390 => x"c348c087",
   391 => x"efc287f8",
   392 => x"c24cbffe",
   393 => x"c25ce7f4",
   394 => x"bf97e3e8",
   395 => x"c231c849",
   396 => x"bf97e2e8",
   397 => x"c249a14a",
   398 => x"bf97e4e8",
   399 => x"7232d04a",
   400 => x"e8c249a1",
   401 => x"4abf97e5",
   402 => x"a17232d8",
   403 => x"9166c449",
   404 => x"bfd3f4c2",
   405 => x"dbf4c281",
   406 => x"ebe8c259",
   407 => x"c84abf97",
   408 => x"eae8c232",
   409 => x"a24bbf97",
   410 => x"ece8c24a",
   411 => x"d04bbf97",
   412 => x"4aa27333",
   413 => x"97ede8c2",
   414 => x"9bcf4bbf",
   415 => x"a27333d8",
   416 => x"dff4c24a",
   417 => x"dbf4c25a",
   418 => x"8ac24abf",
   419 => x"f4c29274",
   420 => x"a17248df",
   421 => x"87cac178",
   422 => x"97d0e8c2",
   423 => x"31c849bf",
   424 => x"97cfe8c2",
   425 => x"49a14abf",
   426 => x"59cef0c2",
   427 => x"bfcaf0c2",
   428 => x"c731c549",
   429 => x"29c981ff",
   430 => x"59e7f4c2",
   431 => x"97d5e8c2",
   432 => x"32c84abf",
   433 => x"97d4e8c2",
   434 => x"4aa24bbf",
   435 => x"6e9266c4",
   436 => x"e3f4c282",
   437 => x"dbf4c25a",
   438 => x"c278c048",
   439 => x"7248d7f4",
   440 => x"f4c278a1",
   441 => x"f4c248e7",
   442 => x"c278bfdb",
   443 => x"c248ebf4",
   444 => x"78bfdff4",
   445 => x"bfc6f0c2",
   446 => x"87c9c002",
   447 => x"30c44874",
   448 => x"c9c07e70",
   449 => x"e3f4c287",
   450 => x"30c448bf",
   451 => x"f0c27e70",
   452 => x"786e48ca",
   453 => x"8ef848c1",
   454 => x"4c264d26",
   455 => x"4f264b26",
   456 => x"5c5b5e0e",
   457 => x"4a710e5d",
   458 => x"bfc6f0c2",
   459 => x"7287cb02",
   460 => x"722bc74b",
   461 => x"9cffc14c",
   462 => x"4b7287c9",
   463 => x"4c722bc8",
   464 => x"c29cffc3",
   465 => x"83bfd3f4",
   466 => x"bfdaf5c0",
   467 => x"87d902ab",
   468 => x"5bdef5c0",
   469 => x"1efee7c2",
   470 => x"fdf04973",
   471 => x"7086c487",
   472 => x"87c50598",
   473 => x"e6c048c0",
   474 => x"c6f0c287",
   475 => x"87d202bf",
   476 => x"91c44974",
   477 => x"81fee7c2",
   478 => x"ffcf4d69",
   479 => x"9dffffff",
   480 => x"497487cb",
   481 => x"e7c291c2",
   482 => x"699f81fe",
   483 => x"fe48754d",
   484 => x"5e0e87c6",
   485 => x"0e5d5c5b",
   486 => x"c04d711e",
   487 => x"cf49c11e",
   488 => x"86c487dc",
   489 => x"029c4c70",
   490 => x"c287c0c1",
   491 => x"754acef0",
   492 => x"87dbe249",
   493 => x"c0029870",
   494 => x"4a7487f1",
   495 => x"4bcb4975",
   496 => x"7087c1e3",
   497 => x"e2c00298",
   498 => x"741ec087",
   499 => x"87c7029c",
   500 => x"c048a6c4",
   501 => x"c487c578",
   502 => x"78c148a6",
   503 => x"ce4966c4",
   504 => x"86c487dc",
   505 => x"059c4c70",
   506 => x"7487c0ff",
   507 => x"e7fc2648",
   508 => x"5b5e0e87",
   509 => x"1e0e5d5c",
   510 => x"059b4b71",
   511 => x"48c087c5",
   512 => x"c887e5c1",
   513 => x"7dc04da3",
   514 => x"c70266d4",
   515 => x"9766d487",
   516 => x"87c505bf",
   517 => x"cfc148c0",
   518 => x"4966d487",
   519 => x"7087f3fd",
   520 => x"c1029c4c",
   521 => x"a4dc87c0",
   522 => x"da7d6949",
   523 => x"a3c449a4",
   524 => x"7a699f4a",
   525 => x"bfc6f0c2",
   526 => x"d487d202",
   527 => x"699f49a4",
   528 => x"ffffc049",
   529 => x"d0487199",
   530 => x"c27e7030",
   531 => x"6e7ec087",
   532 => x"806a4849",
   533 => x"7bc07a70",
   534 => x"6a49a3cc",
   535 => x"49a3d079",
   536 => x"48c179c0",
   537 => x"48c087c2",
   538 => x"87ecfa26",
   539 => x"5c5b5e0e",
   540 => x"4c710e5d",
   541 => x"cac1029c",
   542 => x"49a4c887",
   543 => x"c2c10269",
   544 => x"4a66d087",
   545 => x"d482496c",
   546 => x"66d05aa6",
   547 => x"f0c2b94d",
   548 => x"ff4abfc2",
   549 => x"719972ba",
   550 => x"e4c00299",
   551 => x"4ba4c487",
   552 => x"fbf9496b",
   553 => x"c27b7087",
   554 => x"49bffeef",
   555 => x"7c71816c",
   556 => x"f0c2b975",
   557 => x"ff4abfc2",
   558 => x"719972ba",
   559 => x"dcff0599",
   560 => x"f97c7587",
   561 => x"731e87d2",
   562 => x"9b4b711e",
   563 => x"c887c702",
   564 => x"056949a3",
   565 => x"48c087c5",
   566 => x"c287f7c0",
   567 => x"4abfd7f4",
   568 => x"6949a3c4",
   569 => x"c289c249",
   570 => x"91bffeef",
   571 => x"c24aa271",
   572 => x"49bfc2f0",
   573 => x"a271996b",
   574 => x"def5c04a",
   575 => x"1e66c85a",
   576 => x"d5ea4972",
   577 => x"7086c487",
   578 => x"87c40598",
   579 => x"87c248c0",
   580 => x"c7f848c1",
   581 => x"5b5e0e87",
   582 => x"1e0e5d5c",
   583 => x"66d44b71",
   584 => x"732cc94c",
   585 => x"cfc1029b",
   586 => x"49a3c887",
   587 => x"c7c10269",
   588 => x"4da3d087",
   589 => x"c27d66d4",
   590 => x"49bfc2f0",
   591 => x"4a6bb9ff",
   592 => x"ac717e99",
   593 => x"c087cd03",
   594 => x"a3cc7d7b",
   595 => x"49a3c44a",
   596 => x"87c2796a",
   597 => x"9c748c72",
   598 => x"4987dd02",
   599 => x"fc49731e",
   600 => x"86c487ca",
   601 => x"c74966d4",
   602 => x"cb0299ff",
   603 => x"fee7c287",
   604 => x"fd49731e",
   605 => x"86c487d0",
   606 => x"87dcf626",
   607 => x"5c5b5e0e",
   608 => x"86f00e5d",
   609 => x"c059a6d0",
   610 => x"cc4b66e4",
   611 => x"87ca0266",
   612 => x"7080c848",
   613 => x"05bf6e7e",
   614 => x"48c087c5",
   615 => x"cc87ecc3",
   616 => x"84d04c66",
   617 => x"a6c44973",
   618 => x"c4786c48",
   619 => x"80c48166",
   620 => x"c878bf6e",
   621 => x"c606a966",
   622 => x"66c44987",
   623 => x"c04b7189",
   624 => x"c401abb7",
   625 => x"c2c34887",
   626 => x"4866c487",
   627 => x"7098ffc7",
   628 => x"c1026e7e",
   629 => x"c0c887c9",
   630 => x"71896e49",
   631 => x"fee7c24a",
   632 => x"73856e4d",
   633 => x"c106aab7",
   634 => x"49724a87",
   635 => x"8066c448",
   636 => x"8b727c70",
   637 => x"718ac149",
   638 => x"87d90299",
   639 => x"4866e0c0",
   640 => x"e0c05015",
   641 => x"80c14866",
   642 => x"58a6e4c0",
   643 => x"8ac14972",
   644 => x"e7059971",
   645 => x"d01ec187",
   646 => x"cff94966",
   647 => x"c086c487",
   648 => x"c106abb7",
   649 => x"e0c087e3",
   650 => x"ffc74d66",
   651 => x"c006abb7",
   652 => x"1e7587e2",
   653 => x"fa4966d0",
   654 => x"c0c887cc",
   655 => x"c8486c85",
   656 => x"7c7080c0",
   657 => x"c18bc0c8",
   658 => x"4966d41e",
   659 => x"c887ddf8",
   660 => x"87eec086",
   661 => x"1efee7c2",
   662 => x"f94966d0",
   663 => x"86c487e8",
   664 => x"4afee7c2",
   665 => x"6c484973",
   666 => x"737c7080",
   667 => x"718bc149",
   668 => x"87ce0299",
   669 => x"c17d9712",
   670 => x"c1497385",
   671 => x"0599718b",
   672 => x"b7c087f2",
   673 => x"e1fe01ab",
   674 => x"f048c187",
   675 => x"87c8f28e",
   676 => x"5c5b5e0e",
   677 => x"4b710e5d",
   678 => x"87c7029b",
   679 => x"6d4da3c8",
   680 => x"ff87c505",
   681 => x"87fdc048",
   682 => x"6c4ca3d0",
   683 => x"99ffc749",
   684 => x"6c87d805",
   685 => x"c187c902",
   686 => x"f649731e",
   687 => x"86c487ee",
   688 => x"1efee7c2",
   689 => x"fdf74973",
   690 => x"6c86c487",
   691 => x"04aa6d4a",
   692 => x"48ff87c4",
   693 => x"a2c187cf",
   694 => x"c749727c",
   695 => x"e7c299ff",
   696 => x"699781fe",
   697 => x"87f0f048",
   698 => x"711e731e",
   699 => x"c0029b4b",
   700 => x"f4c287e4",
   701 => x"4a735beb",
   702 => x"efc28ac2",
   703 => x"9249bffe",
   704 => x"bfd7f4c2",
   705 => x"c2807248",
   706 => x"7158eff4",
   707 => x"c230c448",
   708 => x"c058cef0",
   709 => x"f4c287ed",
   710 => x"f4c248e7",
   711 => x"c278bfdb",
   712 => x"c248ebf4",
   713 => x"78bfdff4",
   714 => x"bfc6f0c2",
   715 => x"c287c902",
   716 => x"49bffeef",
   717 => x"87c731c4",
   718 => x"bfe3f4c2",
   719 => x"c231c449",
   720 => x"ef59cef0",
   721 => x"5e0e87d6",
   722 => x"710e5c5b",
   723 => x"724bc04a",
   724 => x"e1c0029a",
   725 => x"49a2da87",
   726 => x"c24b699f",
   727 => x"02bfc6f0",
   728 => x"a2d487cf",
   729 => x"49699f49",
   730 => x"ffffc04c",
   731 => x"c234d09c",
   732 => x"744cc087",
   733 => x"4973b349",
   734 => x"ee87edfd",
   735 => x"5e0e87dc",
   736 => x"0e5d5c5b",
   737 => x"4a7186f4",
   738 => x"9a727ec0",
   739 => x"c287d802",
   740 => x"c048fae7",
   741 => x"f2e7c278",
   742 => x"ebf4c248",
   743 => x"e7c278bf",
   744 => x"f4c248f6",
   745 => x"c278bfe7",
   746 => x"c048dbf0",
   747 => x"caf0c250",
   748 => x"e7c249bf",
   749 => x"714abffa",
   750 => x"cac403aa",
   751 => x"cf497287",
   752 => x"eac00599",
   753 => x"daf5c087",
   754 => x"f2e7c248",
   755 => x"e7c278bf",
   756 => x"e7c21efe",
   757 => x"c249bff2",
   758 => x"c148f2e7",
   759 => x"ff7178a1",
   760 => x"c487f7de",
   761 => x"d6f5c086",
   762 => x"fee7c248",
   763 => x"c087cc78",
   764 => x"48bfd6f5",
   765 => x"c080e0c0",
   766 => x"c258daf5",
   767 => x"48bffae7",
   768 => x"e7c280c1",
   769 => x"562758fe",
   770 => x"bf00000d",
   771 => x"9d4dbf97",
   772 => x"87e3c202",
   773 => x"02ade5c3",
   774 => x"c087dcc2",
   775 => x"4bbfd6f5",
   776 => x"1149a3cb",
   777 => x"05accf4c",
   778 => x"7587d2c1",
   779 => x"c199df49",
   780 => x"c291cd89",
   781 => x"c181cef0",
   782 => x"51124aa3",
   783 => x"124aa3c3",
   784 => x"4aa3c551",
   785 => x"a3c75112",
   786 => x"c951124a",
   787 => x"51124aa3",
   788 => x"124aa3ce",
   789 => x"4aa3d051",
   790 => x"a3d25112",
   791 => x"d451124a",
   792 => x"51124aa3",
   793 => x"124aa3d6",
   794 => x"4aa3d851",
   795 => x"a3dc5112",
   796 => x"de51124a",
   797 => x"51124aa3",
   798 => x"fac07ec1",
   799 => x"c8497487",
   800 => x"ebc00599",
   801 => x"d0497487",
   802 => x"87d10599",
   803 => x"c00266dc",
   804 => x"497387cb",
   805 => x"700f66dc",
   806 => x"d3c00298",
   807 => x"c0056e87",
   808 => x"f0c287c6",
   809 => x"50c048ce",
   810 => x"bfd6f5c0",
   811 => x"87e1c248",
   812 => x"48dbf0c2",
   813 => x"c27e50c0",
   814 => x"49bfcaf0",
   815 => x"bffae7c2",
   816 => x"04aa714a",
   817 => x"c287f6fb",
   818 => x"05bfebf4",
   819 => x"c287c8c0",
   820 => x"02bfc6f0",
   821 => x"c287f8c1",
   822 => x"49bff6e7",
   823 => x"7087c1e9",
   824 => x"fae7c249",
   825 => x"48a6c459",
   826 => x"bff6e7c2",
   827 => x"c6f0c278",
   828 => x"d8c002bf",
   829 => x"4966c487",
   830 => x"ffffffcf",
   831 => x"02a999f8",
   832 => x"c087c5c0",
   833 => x"87e1c04c",
   834 => x"dcc04cc1",
   835 => x"4966c487",
   836 => x"99f8ffcf",
   837 => x"c8c002a9",
   838 => x"48a6c887",
   839 => x"c5c078c0",
   840 => x"48a6c887",
   841 => x"66c878c1",
   842 => x"059c744c",
   843 => x"c487e0c0",
   844 => x"89c24966",
   845 => x"bffeefc2",
   846 => x"f4c2914a",
   847 => x"c24abfd7",
   848 => x"7248f2e7",
   849 => x"e7c278a1",
   850 => x"78c048fa",
   851 => x"c087def9",
   852 => x"e78ef448",
   853 => x"000087c2",
   854 => x"ffff0000",
   855 => x"0d66ffff",
   856 => x"0d6f0000",
   857 => x"41460000",
   858 => x"20323354",
   859 => x"46002020",
   860 => x"36315441",
   861 => x"00202020",
   862 => x"f0f4c21e",
   863 => x"a8dd48bf",
   864 => x"c187c905",
   865 => x"7087e3c2",
   866 => x"87c84a49",
   867 => x"c348d4ff",
   868 => x"4a6878ff",
   869 => x"4f264872",
   870 => x"f0f4c21e",
   871 => x"a8dd48bf",
   872 => x"c187c605",
   873 => x"d987efc1",
   874 => x"48d4ff87",
   875 => x"ff78ffc3",
   876 => x"e1c048d0",
   877 => x"48d4ff78",
   878 => x"f4c278d4",
   879 => x"d4ff48ef",
   880 => x"4f2650bf",
   881 => x"48d0ff1e",
   882 => x"2678e0c0",
   883 => x"e7fe1e4f",
   884 => x"99497087",
   885 => x"c087c602",
   886 => x"f105a9fb",
   887 => x"26487187",
   888 => x"5b5e0e4f",
   889 => x"4b710e5c",
   890 => x"cbfe4cc0",
   891 => x"99497087",
   892 => x"87f9c002",
   893 => x"02a9ecc0",
   894 => x"c087f2c0",
   895 => x"c002a9fb",
   896 => x"66cc87eb",
   897 => x"c703acb7",
   898 => x"0266d087",
   899 => x"537187c2",
   900 => x"c2029971",
   901 => x"fd84c187",
   902 => x"497087de",
   903 => x"87cd0299",
   904 => x"02a9ecc0",
   905 => x"fbc087c7",
   906 => x"d5ff05a9",
   907 => x"0266d087",
   908 => x"97c087c3",
   909 => x"a9ecc07b",
   910 => x"7487c405",
   911 => x"7487c54a",
   912 => x"8a0ac04a",
   913 => x"87c24872",
   914 => x"4c264d26",
   915 => x"4f264b26",
   916 => x"87e4fc1e",
   917 => x"f0c04970",
   918 => x"ca04a9b7",
   919 => x"b7f9c087",
   920 => x"87c301a9",
   921 => x"c189f0c0",
   922 => x"04a9b7c1",
   923 => x"dac187ca",
   924 => x"c301a9b7",
   925 => x"89f7c087",
   926 => x"4f264871",
   927 => x"5c5b5e0e",
   928 => x"fc4c710e",
   929 => x"1ec187d2",
   930 => x"741e66d0",
   931 => x"87d1fd49",
   932 => x"4b7086c8",
   933 => x"c087edfc",
   934 => x"c203abb7",
   935 => x"cc8b0b87",
   936 => x"03abb766",
   937 => x"a37487cf",
   938 => x"c083c149",
   939 => x"66cc51e0",
   940 => x"f104abb7",
   941 => x"49a37487",
   942 => x"cdfe51c0",
   943 => x"5b5e0e87",
   944 => x"4a710e5c",
   945 => x"724cd4ff",
   946 => x"87e9c049",
   947 => x"029b4b70",
   948 => x"8bc187c2",
   949 => x"c548d0ff",
   950 => x"7cd5c178",
   951 => x"31c64973",
   952 => x"97d7e7c1",
   953 => x"71484abf",
   954 => x"ff7c70b0",
   955 => x"78c448d0",
   956 => x"d5fd4873",
   957 => x"5b5e0e87",
   958 => x"f40e5d5c",
   959 => x"c44c7186",
   960 => x"78c048a6",
   961 => x"6e7ea4c8",
   962 => x"c149bf97",
   963 => x"dd05a9c1",
   964 => x"49a4c987",
   965 => x"c1496997",
   966 => x"d105a9d2",
   967 => x"49a4ca87",
   968 => x"c1496997",
   969 => x"c505a9c3",
   970 => x"c248df87",
   971 => x"e7f987e1",
   972 => x"c04bc087",
   973 => x"bf97d4ff",
   974 => x"04a9c049",
   975 => x"ccfa87cf",
   976 => x"c083c187",
   977 => x"bf97d4ff",
   978 => x"f106ab49",
   979 => x"d4ffc087",
   980 => x"cf02bf97",
   981 => x"87e0f887",
   982 => x"02994970",
   983 => x"ecc087c6",
   984 => x"87f105a9",
   985 => x"cff84bc0",
   986 => x"f84d7087",
   987 => x"a6cc87ca",
   988 => x"87c4f858",
   989 => x"83c14a70",
   990 => x"49bf976e",
   991 => x"87c702ad",
   992 => x"05adffc0",
   993 => x"c987eac0",
   994 => x"699749a4",
   995 => x"a966c849",
   996 => x"4887c702",
   997 => x"05a8ffc0",
   998 => x"a4ca87d7",
   999 => x"49699749",
  1000 => x"87c602aa",
  1001 => x"05aaffc0",
  1002 => x"a6c487c7",
  1003 => x"d378c148",
  1004 => x"adecc087",
  1005 => x"c087c602",
  1006 => x"c705adfb",
  1007 => x"c44bc087",
  1008 => x"78c148a6",
  1009 => x"fe0266c4",
  1010 => x"f7f787dc",
  1011 => x"f4487387",
  1012 => x"87f4f98e",
  1013 => x"5b5e0e00",
  1014 => x"1e0e5d5c",
  1015 => x"d4ff4d71",
  1016 => x"c21e754b",
  1017 => x"e049f4f4",
  1018 => x"86c487c7",
  1019 => x"c4029870",
  1020 => x"f4c287c8",
  1021 => x"754cbffc",
  1022 => x"87c1fb49",
  1023 => x"c005a8de",
  1024 => x"497587eb",
  1025 => x"87c0f6c0",
  1026 => x"db029870",
  1027 => x"d8f9c287",
  1028 => x"e1c01ebf",
  1029 => x"cff3c049",
  1030 => x"c186c487",
  1031 => x"c048d7e7",
  1032 => x"e4f9c250",
  1033 => x"87edfe49",
  1034 => x"cfc348c1",
  1035 => x"48d0ff87",
  1036 => x"d6c178c5",
  1037 => x"754ac07b",
  1038 => x"7b1149a2",
  1039 => x"b7cb82c1",
  1040 => x"87f304aa",
  1041 => x"ffc34acc",
  1042 => x"c082c17b",
  1043 => x"04aab7e0",
  1044 => x"d0ff87f4",
  1045 => x"c378c448",
  1046 => x"78c57bff",
  1047 => x"c17bd3c1",
  1048 => x"7478c47b",
  1049 => x"c0c2029c",
  1050 => x"fee7c287",
  1051 => x"4dc0c87e",
  1052 => x"acb7c08c",
  1053 => x"c887c603",
  1054 => x"c04da4c0",
  1055 => x"adc0c84c",
  1056 => x"c287dc05",
  1057 => x"bf97eff4",
  1058 => x"0299d049",
  1059 => x"1ec087d1",
  1060 => x"49f4f4c2",
  1061 => x"c487efe0",
  1062 => x"4a497086",
  1063 => x"c287eec0",
  1064 => x"c21efee7",
  1065 => x"e049f4f4",
  1066 => x"86c487dc",
  1067 => x"ff4a4970",
  1068 => x"c5c848d0",
  1069 => x"7bd4c178",
  1070 => x"7bbf976e",
  1071 => x"80c1486e",
  1072 => x"8dc17e70",
  1073 => x"87f0ff05",
  1074 => x"c448d0ff",
  1075 => x"059a7278",
  1076 => x"48c087c5",
  1077 => x"c187e5c0",
  1078 => x"f4f4c21e",
  1079 => x"cbdeff49",
  1080 => x"7486c487",
  1081 => x"c0fe059c",
  1082 => x"48d0ff87",
  1083 => x"d3c178c5",
  1084 => x"c47bc07b",
  1085 => x"c048c178",
  1086 => x"48c087c2",
  1087 => x"264d2626",
  1088 => x"264b264c",
  1089 => x"5b5e0e4f",
  1090 => x"1e0e5d5c",
  1091 => x"4cc04b71",
  1092 => x"c004ab4d",
  1093 => x"fbc087e8",
  1094 => x"9d751ef5",
  1095 => x"c087c402",
  1096 => x"c187c24a",
  1097 => x"e949724a",
  1098 => x"86c487d4",
  1099 => x"84c17e70",
  1100 => x"87c2056e",
  1101 => x"85c14c73",
  1102 => x"ff06ac73",
  1103 => x"486e87d8",
  1104 => x"87f9fe26",
  1105 => x"c44a711e",
  1106 => x"87c50566",
  1107 => x"c4fa4972",
  1108 => x"0e4f2687",
  1109 => x"5d5c5b5e",
  1110 => x"4c711e0e",
  1111 => x"c291de49",
  1112 => x"714ddcf5",
  1113 => x"026d9785",
  1114 => x"c287dcc1",
  1115 => x"4abfc8f5",
  1116 => x"49728274",
  1117 => x"7087cefe",
  1118 => x"c0026e7e",
  1119 => x"f5c287f2",
  1120 => x"4a6e4bd0",
  1121 => x"fcfe49cb",
  1122 => x"4b7487de",
  1123 => x"e7c193cb",
  1124 => x"83c483e7",
  1125 => x"7bcbc7c1",
  1126 => x"cbc14974",
  1127 => x"7b7587d7",
  1128 => x"97d8e7c1",
  1129 => x"c21e49bf",
  1130 => x"fe49d0f5",
  1131 => x"86c487d6",
  1132 => x"cac14974",
  1133 => x"49c087ff",
  1134 => x"87deccc1",
  1135 => x"48f0f4c2",
  1136 => x"49c178c0",
  1137 => x"2687cfdd",
  1138 => x"4c87f2fc",
  1139 => x"6964616f",
  1140 => x"2e2e676e",
  1141 => x"5e0e002e",
  1142 => x"710e5c5b",
  1143 => x"f5c24a4b",
  1144 => x"7282bfc8",
  1145 => x"87ddfc49",
  1146 => x"029c4c70",
  1147 => x"e54987c4",
  1148 => x"f5c287d4",
  1149 => x"78c048c8",
  1150 => x"d9dc49c1",
  1151 => x"87fffb87",
  1152 => x"5c5b5e0e",
  1153 => x"86f40e5d",
  1154 => x"4dfee7c2",
  1155 => x"a6c44cc0",
  1156 => x"c278c048",
  1157 => x"49bfc8f5",
  1158 => x"c106a9c0",
  1159 => x"e7c287c1",
  1160 => x"029848fe",
  1161 => x"c087f8c0",
  1162 => x"c81ef5fb",
  1163 => x"87c70266",
  1164 => x"c048a6c4",
  1165 => x"c487c578",
  1166 => x"78c148a6",
  1167 => x"e44966c4",
  1168 => x"86c487fc",
  1169 => x"84c14d70",
  1170 => x"c14866c4",
  1171 => x"58a6c880",
  1172 => x"bfc8f5c2",
  1173 => x"c603ac49",
  1174 => x"059d7587",
  1175 => x"c087c8ff",
  1176 => x"029d754c",
  1177 => x"c087e0c3",
  1178 => x"c81ef5fb",
  1179 => x"87c70266",
  1180 => x"c048a6cc",
  1181 => x"cc87c578",
  1182 => x"78c148a6",
  1183 => x"e34966cc",
  1184 => x"86c487fc",
  1185 => x"026e7e70",
  1186 => x"6e87e9c2",
  1187 => x"9781cb49",
  1188 => x"99d04969",
  1189 => x"87d6c102",
  1190 => x"4ad6c7c1",
  1191 => x"91cb4974",
  1192 => x"81e7e7c1",
  1193 => x"81c87972",
  1194 => x"7451ffc3",
  1195 => x"c291de49",
  1196 => x"714ddcf5",
  1197 => x"97c1c285",
  1198 => x"49a5c17d",
  1199 => x"c251e0c0",
  1200 => x"bf97cef0",
  1201 => x"c187d202",
  1202 => x"4ba5c284",
  1203 => x"4acef0c2",
  1204 => x"f7fe49db",
  1205 => x"dbc187d2",
  1206 => x"49a5cd87",
  1207 => x"84c151c0",
  1208 => x"6e4ba5c2",
  1209 => x"fe49cb4a",
  1210 => x"c187fdf6",
  1211 => x"c5c187c6",
  1212 => x"49744ad3",
  1213 => x"e7c191cb",
  1214 => x"797281e7",
  1215 => x"97cef0c2",
  1216 => x"87d802bf",
  1217 => x"91de4974",
  1218 => x"f5c284c1",
  1219 => x"83714bdc",
  1220 => x"4acef0c2",
  1221 => x"f6fe49dd",
  1222 => x"87d887ce",
  1223 => x"93de4b74",
  1224 => x"83dcf5c2",
  1225 => x"c049a3cb",
  1226 => x"7384c151",
  1227 => x"49cb4a6e",
  1228 => x"87f4f5fe",
  1229 => x"c14866c4",
  1230 => x"58a6c880",
  1231 => x"c003acc7",
  1232 => x"056e87c5",
  1233 => x"7487e0fc",
  1234 => x"f68ef448",
  1235 => x"731e87ef",
  1236 => x"494b711e",
  1237 => x"e7c191cb",
  1238 => x"a1c881e7",
  1239 => x"d7e7c14a",
  1240 => x"c9501248",
  1241 => x"ffc04aa1",
  1242 => x"501248d4",
  1243 => x"e7c181ca",
  1244 => x"501148d8",
  1245 => x"97d8e7c1",
  1246 => x"c01e49bf",
  1247 => x"87c4f749",
  1248 => x"48f0f4c2",
  1249 => x"49c178de",
  1250 => x"2687cbd6",
  1251 => x"1e87f2f5",
  1252 => x"cb494a71",
  1253 => x"e7e7c191",
  1254 => x"1181c881",
  1255 => x"f4f4c248",
  1256 => x"c8f5c258",
  1257 => x"c178c048",
  1258 => x"87ead549",
  1259 => x"c01e4f26",
  1260 => x"e5c4c149",
  1261 => x"1e4f2687",
  1262 => x"d2029971",
  1263 => x"fce8c187",
  1264 => x"f750c048",
  1265 => x"cfcec180",
  1266 => x"e0e7c140",
  1267 => x"c187ce78",
  1268 => x"c148f8e8",
  1269 => x"fc78d9e7",
  1270 => x"eecec180",
  1271 => x"0e4f2678",
  1272 => x"0e5c5b5e",
  1273 => x"cb4a4c71",
  1274 => x"e7e7c192",
  1275 => x"49a2c882",
  1276 => x"974ba2c9",
  1277 => x"971e4b6b",
  1278 => x"ca1e4969",
  1279 => x"c0491282",
  1280 => x"c087c5e5",
  1281 => x"87ced449",
  1282 => x"c1c14974",
  1283 => x"8ef887e7",
  1284 => x"1e87ecf3",
  1285 => x"4b711e73",
  1286 => x"87c3ff49",
  1287 => x"fefe4973",
  1288 => x"87ddf387",
  1289 => x"711e731e",
  1290 => x"4aa3c64b",
  1291 => x"c187db02",
  1292 => x"87d6028a",
  1293 => x"dac1028a",
  1294 => x"c0028a87",
  1295 => x"028a87fc",
  1296 => x"8a87e1c0",
  1297 => x"c187cb02",
  1298 => x"49c787db",
  1299 => x"c187c0fd",
  1300 => x"f5c287de",
  1301 => x"c102bfc8",
  1302 => x"c14887cb",
  1303 => x"ccf5c288",
  1304 => x"87c1c158",
  1305 => x"bfccf5c2",
  1306 => x"87f9c002",
  1307 => x"bfc8f5c2",
  1308 => x"c280c148",
  1309 => x"c058ccf5",
  1310 => x"f5c287eb",
  1311 => x"c649bfc8",
  1312 => x"ccf5c289",
  1313 => x"a9b7c059",
  1314 => x"c287da03",
  1315 => x"c048c8f5",
  1316 => x"c287d278",
  1317 => x"02bfccf5",
  1318 => x"f5c287cb",
  1319 => x"c648bfc8",
  1320 => x"ccf5c280",
  1321 => x"d149c058",
  1322 => x"497387ec",
  1323 => x"87c5ffc0",
  1324 => x"1e87cef1",
  1325 => x"4b711e73",
  1326 => x"48f0f4c2",
  1327 => x"49c078dd",
  1328 => x"7387d3d1",
  1329 => x"ecfec049",
  1330 => x"87f5f087",
  1331 => x"5c5b5e0e",
  1332 => x"cc4c710e",
  1333 => x"4b741e66",
  1334 => x"e7c193cb",
  1335 => x"a3c483e7",
  1336 => x"fe496a4a",
  1337 => x"c187d1ef",
  1338 => x"c87bcecd",
  1339 => x"66d449a3",
  1340 => x"49a3c951",
  1341 => x"ca5166d8",
  1342 => x"66dc49a3",
  1343 => x"feef2651",
  1344 => x"5b5e0e87",
  1345 => x"ff0e5d5c",
  1346 => x"a6dc86cc",
  1347 => x"48a6c859",
  1348 => x"80c478c0",
  1349 => x"7866c8c1",
  1350 => x"78c180c4",
  1351 => x"78c180c4",
  1352 => x"48ccf5c2",
  1353 => x"f4c278c1",
  1354 => x"de48bff0",
  1355 => x"87cb05a8",
  1356 => x"7087cdf3",
  1357 => x"59a6cc49",
  1358 => x"e187d6ce",
  1359 => x"cce287da",
  1360 => x"87f4e087",
  1361 => x"fbc04c70",
  1362 => x"d8c102ac",
  1363 => x"0566d887",
  1364 => x"c087cac1",
  1365 => x"1ec11e1e",
  1366 => x"1ecae9c1",
  1367 => x"ebfd49c0",
  1368 => x"c086d087",
  1369 => x"d902acfb",
  1370 => x"66c4c187",
  1371 => x"6a82c44a",
  1372 => x"7481c749",
  1373 => x"d81ec151",
  1374 => x"c8496a1e",
  1375 => x"87e1e181",
  1376 => x"c8c186c8",
  1377 => x"a8c04866",
  1378 => x"c887c701",
  1379 => x"78c148a6",
  1380 => x"c8c187ce",
  1381 => x"88c14866",
  1382 => x"c358a6d0",
  1383 => x"87ede087",
  1384 => x"c248a6d0",
  1385 => x"029c7478",
  1386 => x"c887e2cc",
  1387 => x"ccc14866",
  1388 => x"cc03a866",
  1389 => x"a6c487d7",
  1390 => x"d878c048",
  1391 => x"ff78c080",
  1392 => x"7087f5de",
  1393 => x"4866d84c",
  1394 => x"c605a8dd",
  1395 => x"48a6dc87",
  1396 => x"c17866d8",
  1397 => x"c005acd0",
  1398 => x"deff87eb",
  1399 => x"deff87da",
  1400 => x"4c7087d6",
  1401 => x"05acecc0",
  1402 => x"dfff87c6",
  1403 => x"4c7087df",
  1404 => x"05acd0c1",
  1405 => x"66d487c8",
  1406 => x"d880c148",
  1407 => x"d0c158a6",
  1408 => x"d5ff02ac",
  1409 => x"a6e0c087",
  1410 => x"7866d848",
  1411 => x"c04866dc",
  1412 => x"05a866e0",
  1413 => x"c087c8ca",
  1414 => x"c048a6e4",
  1415 => x"c080c478",
  1416 => x"c04d7478",
  1417 => x"c9028dfb",
  1418 => x"8dc987ce",
  1419 => x"c287db02",
  1420 => x"f7c1028d",
  1421 => x"028dc987",
  1422 => x"c487d1c4",
  1423 => x"c2c1028d",
  1424 => x"028dc187",
  1425 => x"c887c5c4",
  1426 => x"66c887e8",
  1427 => x"c191cb49",
  1428 => x"c48166c4",
  1429 => x"7e6a4aa1",
  1430 => x"e4c11e71",
  1431 => x"66c448c9",
  1432 => x"4aa1cc49",
  1433 => x"aa714120",
  1434 => x"87f8ff05",
  1435 => x"49265110",
  1436 => x"79f3d2c1",
  1437 => x"87d5ddff",
  1438 => x"e8c04c70",
  1439 => x"78c148a6",
  1440 => x"c487f5c7",
  1441 => x"f0c048a6",
  1442 => x"ebdbff78",
  1443 => x"c04c7087",
  1444 => x"c002acec",
  1445 => x"a6c887c3",
  1446 => x"acecc05c",
  1447 => x"ff87cd02",
  1448 => x"7087d5db",
  1449 => x"acecc04c",
  1450 => x"87f3ff05",
  1451 => x"02acecc0",
  1452 => x"ff87c4c0",
  1453 => x"c487c1db",
  1454 => x"66d81e66",
  1455 => x"66d81e49",
  1456 => x"e9c11e49",
  1457 => x"66d81eca",
  1458 => x"87c0f849",
  1459 => x"1eca1ec0",
  1460 => x"4966e0c0",
  1461 => x"dcc191cb",
  1462 => x"a6d88166",
  1463 => x"78a1c448",
  1464 => x"49bf66d8",
  1465 => x"87f9dbff",
  1466 => x"b7c086d8",
  1467 => x"cbc106a8",
  1468 => x"de1ec187",
  1469 => x"bf66c81e",
  1470 => x"e4dbff49",
  1471 => x"7086c887",
  1472 => x"08c04849",
  1473 => x"a6ecc088",
  1474 => x"a8b7c058",
  1475 => x"87ecc006",
  1476 => x"4866e8c0",
  1477 => x"03a8b7dd",
  1478 => x"6e87e1c0",
  1479 => x"e8c049bf",
  1480 => x"e0c08166",
  1481 => x"66e8c051",
  1482 => x"6e81c149",
  1483 => x"c1c281bf",
  1484 => x"66e8c051",
  1485 => x"6e81c249",
  1486 => x"51c081bf",
  1487 => x"c14866d0",
  1488 => x"58a6d480",
  1489 => x"c180d848",
  1490 => x"87ecc478",
  1491 => x"87c0dcff",
  1492 => x"58a6ecc0",
  1493 => x"87f8dbff",
  1494 => x"58a6f0c0",
  1495 => x"05a8ecc0",
  1496 => x"a687c9c0",
  1497 => x"66e8c048",
  1498 => x"87c4c078",
  1499 => x"87c8d8ff",
  1500 => x"cb4966c8",
  1501 => x"66c4c191",
  1502 => x"c8807148",
  1503 => x"66c458a6",
  1504 => x"c482c84a",
  1505 => x"81ca4966",
  1506 => x"5166e8c0",
  1507 => x"4966ecc0",
  1508 => x"e8c081c1",
  1509 => x"48c18966",
  1510 => x"49703071",
  1511 => x"977189c1",
  1512 => x"f8f8c27a",
  1513 => x"e8c049bf",
  1514 => x"6a972966",
  1515 => x"9871484a",
  1516 => x"58a6f4c0",
  1517 => x"c44966c4",
  1518 => x"c07e6981",
  1519 => x"dc4866e0",
  1520 => x"c002a866",
  1521 => x"a6dc87c8",
  1522 => x"c078c048",
  1523 => x"a6dc87c5",
  1524 => x"dc78c148",
  1525 => x"e0c01e66",
  1526 => x"4966c81e",
  1527 => x"87c1d8ff",
  1528 => x"4c7086c8",
  1529 => x"06acb7c0",
  1530 => x"6e87d6c1",
  1531 => x"70807448",
  1532 => x"49e0c07e",
  1533 => x"4b6e8974",
  1534 => x"4ac6e4c1",
  1535 => x"e7e2fe71",
  1536 => x"c2486e87",
  1537 => x"c07e7080",
  1538 => x"c14866e4",
  1539 => x"a6e8c080",
  1540 => x"66f0c058",
  1541 => x"7081c149",
  1542 => x"c5c002a9",
  1543 => x"c04dc087",
  1544 => x"4dc187c2",
  1545 => x"a4c21e75",
  1546 => x"48e0c049",
  1547 => x"49708871",
  1548 => x"4966c81e",
  1549 => x"87e9d6ff",
  1550 => x"b7c086c8",
  1551 => x"c6ff01a8",
  1552 => x"66e4c087",
  1553 => x"87d3c002",
  1554 => x"c94966c4",
  1555 => x"66e4c081",
  1556 => x"4866c451",
  1557 => x"78dfcfc1",
  1558 => x"c487cec0",
  1559 => x"81c94966",
  1560 => x"66c451c2",
  1561 => x"d3d0c148",
  1562 => x"a6e8c078",
  1563 => x"c078c148",
  1564 => x"d5ff87c6",
  1565 => x"4c7087d7",
  1566 => x"0266e8c0",
  1567 => x"c887f5c0",
  1568 => x"66cc4866",
  1569 => x"cbc004a8",
  1570 => x"4866c887",
  1571 => x"a6cc80c1",
  1572 => x"87e0c058",
  1573 => x"c14866cc",
  1574 => x"58a6d088",
  1575 => x"c187d5c0",
  1576 => x"c005acc6",
  1577 => x"66d087c8",
  1578 => x"d480c148",
  1579 => x"d4ff58a6",
  1580 => x"4c7087db",
  1581 => x"c14866d4",
  1582 => x"58a6d880",
  1583 => x"c0029c74",
  1584 => x"66c887cb",
  1585 => x"66ccc148",
  1586 => x"e9f304a8",
  1587 => x"f3d3ff87",
  1588 => x"4866c887",
  1589 => x"c003a8c7",
  1590 => x"f5c287e5",
  1591 => x"78c048cc",
  1592 => x"cb4966c8",
  1593 => x"66c4c191",
  1594 => x"4aa1c481",
  1595 => x"52c04a6a",
  1596 => x"4866c879",
  1597 => x"a6cc80c1",
  1598 => x"04a8c758",
  1599 => x"ff87dbff",
  1600 => x"dfff8ecc",
  1601 => x"203a87f7",
  1602 => x"50494400",
  1603 => x"69775320",
  1604 => x"65686374",
  1605 => x"731e0073",
  1606 => x"9b4b711e",
  1607 => x"c287c602",
  1608 => x"c048c8f5",
  1609 => x"c21ec778",
  1610 => x"49bfc8f5",
  1611 => x"e7e7c11e",
  1612 => x"f0f4c21e",
  1613 => x"c8ef49bf",
  1614 => x"c286cc87",
  1615 => x"49bff0f4",
  1616 => x"7387f4e9",
  1617 => x"87c8029b",
  1618 => x"49e7e7c1",
  1619 => x"87f7edc0",
  1620 => x"87eddeff",
  1621 => x"87d1c71e",
  1622 => x"f9fe49c1",
  1623 => x"e2e5fe87",
  1624 => x"02987087",
  1625 => x"ecfe87cd",
  1626 => x"987087fb",
  1627 => x"c187c402",
  1628 => x"c087c24a",
  1629 => x"059a724a",
  1630 => x"1ec087ce",
  1631 => x"49e9e6c1",
  1632 => x"87e1f9c0",
  1633 => x"87fe86c4",
  1634 => x"87c4fcc0",
  1635 => x"e6c11ec0",
  1636 => x"f9c049f4",
  1637 => x"1ec087cf",
  1638 => x"87cafec0",
  1639 => x"f9c04970",
  1640 => x"c3c387c3",
  1641 => x"268ef887",
  1642 => x"2044534f",
  1643 => x"6c696166",
  1644 => x"002e6465",
  1645 => x"746f6f42",
  1646 => x"2e676e69",
  1647 => x"1e002e2e",
  1648 => x"48c8f5c2",
  1649 => x"f4c278c0",
  1650 => x"78c048f0",
  1651 => x"c087c5fe",
  1652 => x"c087f1ff",
  1653 => x"004f2648",
  1654 => x"45208000",
  1655 => x"00746978",
  1656 => x"61422080",
  1657 => x"8f006b63",
  1658 => x"5c000013",
  1659 => x"0000002d",
  1660 => x"138f0000",
  1661 => x"2d7a0000",
  1662 => x"00000000",
  1663 => x"00138f00",
  1664 => x"002d9800",
  1665 => x"00000000",
  1666 => x"0000138f",
  1667 => x"00002db6",
  1668 => x"8f000000",
  1669 => x"d4000013",
  1670 => x"0000002d",
  1671 => x"138f0000",
  1672 => x"2df20000",
  1673 => x"00000000",
  1674 => x"00138f00",
  1675 => x"002e1000",
  1676 => x"00000000",
  1677 => x"0000138f",
  1678 => x"00000000",
  1679 => x"24000000",
  1680 => x"00000014",
  1681 => x"00000000",
  1682 => x"6f4c0000",
  1683 => x"2a206461",
  1684 => x"fe1e002e",
  1685 => x"78c048f0",
  1686 => x"097909cd",
  1687 => x"1e1e4f26",
  1688 => x"7ebff0fe",
  1689 => x"4f262648",
  1690 => x"48f0fe1e",
  1691 => x"4f2678c1",
  1692 => x"48f0fe1e",
  1693 => x"4f2678c0",
  1694 => x"c04a711e",
  1695 => x"4f265252",
  1696 => x"5c5b5e0e",
  1697 => x"86f40e5d",
  1698 => x"6d974d71",
  1699 => x"4ca5c17e",
  1700 => x"c8486c97",
  1701 => x"486e58a6",
  1702 => x"05a866c4",
  1703 => x"48ff87c5",
  1704 => x"ff87e6c0",
  1705 => x"a5c287ca",
  1706 => x"4b6c9749",
  1707 => x"974ba371",
  1708 => x"6c974b6b",
  1709 => x"c1486e7e",
  1710 => x"58a6c880",
  1711 => x"a6cc98c7",
  1712 => x"7c977058",
  1713 => x"7387e1fe",
  1714 => x"268ef448",
  1715 => x"264c264d",
  1716 => x"0e4f264b",
  1717 => x"0e5c5b5e",
  1718 => x"4c7186f4",
  1719 => x"c34a66d8",
  1720 => x"a4c29aff",
  1721 => x"496c974b",
  1722 => x"7249a173",
  1723 => x"7e6c9751",
  1724 => x"80c1486e",
  1725 => x"c758a6c8",
  1726 => x"58a6cc98",
  1727 => x"8ef45470",
  1728 => x"1e87caff",
  1729 => x"87e8fd1e",
  1730 => x"494abfe0",
  1731 => x"99c0e0c0",
  1732 => x"7287cb02",
  1733 => x"eef8c21e",
  1734 => x"87f7fe49",
  1735 => x"fdfc86c4",
  1736 => x"fd7e7087",
  1737 => x"262687c2",
  1738 => x"f8c21e4f",
  1739 => x"c7fd49ee",
  1740 => x"c3ecc187",
  1741 => x"87dafc49",
  1742 => x"2687c8c4",
  1743 => x"d0ff1e4f",
  1744 => x"78e1c848",
  1745 => x"c548d4ff",
  1746 => x"0266c478",
  1747 => x"e0c387c3",
  1748 => x"0266c878",
  1749 => x"d4ff87c6",
  1750 => x"78f0c348",
  1751 => x"7148d4ff",
  1752 => x"48d0ff78",
  1753 => x"c078e1c8",
  1754 => x"4f2678e0",
  1755 => x"5c5b5e0e",
  1756 => x"c24c710e",
  1757 => x"fc49eef8",
  1758 => x"4a7087c6",
  1759 => x"04aab7c0",
  1760 => x"c387e3c2",
  1761 => x"c905aae0",
  1762 => x"f6f0c187",
  1763 => x"c278c148",
  1764 => x"f0c387d4",
  1765 => x"87c905aa",
  1766 => x"48f2f0c1",
  1767 => x"f5c178c1",
  1768 => x"f6f0c187",
  1769 => x"87c702bf",
  1770 => x"c0c24b72",
  1771 => x"7287c2b3",
  1772 => x"059c744b",
  1773 => x"f0c187d1",
  1774 => x"c11ebff2",
  1775 => x"1ebff6f0",
  1776 => x"f8fd4972",
  1777 => x"c186c887",
  1778 => x"02bff2f0",
  1779 => x"7387e0c0",
  1780 => x"29b7c449",
  1781 => x"d2f2c191",
  1782 => x"cf4a7381",
  1783 => x"c192c29a",
  1784 => x"70307248",
  1785 => x"72baff4a",
  1786 => x"70986948",
  1787 => x"7387db79",
  1788 => x"29b7c449",
  1789 => x"d2f2c191",
  1790 => x"cf4a7381",
  1791 => x"c392c29a",
  1792 => x"70307248",
  1793 => x"b069484a",
  1794 => x"f0c17970",
  1795 => x"78c048f6",
  1796 => x"48f2f0c1",
  1797 => x"f8c278c0",
  1798 => x"e3f949ee",
  1799 => x"c04a7087",
  1800 => x"fd03aab7",
  1801 => x"48c087dd",
  1802 => x"4d2687c2",
  1803 => x"4b264c26",
  1804 => x"00004f26",
  1805 => x"00000000",
  1806 => x"711e0000",
  1807 => x"ebfc494a",
  1808 => x"1e4f2687",
  1809 => x"49724ac0",
  1810 => x"f2c191c4",
  1811 => x"79c081d2",
  1812 => x"b7d082c1",
  1813 => x"87ee04aa",
  1814 => x"5e0e4f26",
  1815 => x"0e5d5c5b",
  1816 => x"cbf84d71",
  1817 => x"c44a7587",
  1818 => x"c1922ab7",
  1819 => x"7582d2f2",
  1820 => x"c29ccf4c",
  1821 => x"4b496a94",
  1822 => x"9bc32b74",
  1823 => x"307448c2",
  1824 => x"bcff4c70",
  1825 => x"98714874",
  1826 => x"dbf77a70",
  1827 => x"fe487387",
  1828 => x"000087d8",
  1829 => x"00000000",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00000000",
  1834 => x"00000000",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"00000000",
  1842 => x"00000000",
  1843 => x"00000000",
  1844 => x"ff1e0000",
  1845 => x"e1c848d0",
  1846 => x"ff487178",
  1847 => x"c47808d4",
  1848 => x"d4ff4866",
  1849 => x"4f267808",
  1850 => x"c44a711e",
  1851 => x"721e4966",
  1852 => x"87deff49",
  1853 => x"c048d0ff",
  1854 => x"262678e0",
  1855 => x"1e731e4f",
  1856 => x"66c84b71",
  1857 => x"4a731e49",
  1858 => x"49a2e0c1",
  1859 => x"2687d9ff",
  1860 => x"4d2687c4",
  1861 => x"4b264c26",
  1862 => x"ff1e4f26",
  1863 => x"ffc34ad4",
  1864 => x"48d0ff7a",
  1865 => x"de78e1c0",
  1866 => x"f8f8c27a",
  1867 => x"48497abf",
  1868 => x"7a7028c8",
  1869 => x"28d04871",
  1870 => x"48717a70",
  1871 => x"7a7028d8",
  1872 => x"c048d0ff",
  1873 => x"4f2678e0",
  1874 => x"5c5b5e0e",
  1875 => x"4c710e5d",
  1876 => x"bff8f8c2",
  1877 => x"2b744b4d",
  1878 => x"c19b66d0",
  1879 => x"ab66d483",
  1880 => x"c087c204",
  1881 => x"d04a744b",
  1882 => x"31724966",
  1883 => x"9975b9ff",
  1884 => x"30724873",
  1885 => x"71484a70",
  1886 => x"fcf8c2b0",
  1887 => x"87dafe58",
  1888 => x"4c264d26",
  1889 => x"4f264b26",
  1890 => x"5c5b5e0e",
  1891 => x"711e0e5d",
  1892 => x"fcf8c24c",
  1893 => x"c04ac04b",
  1894 => x"ccfe49f4",
  1895 => x"1e7487e7",
  1896 => x"49fcf8c2",
  1897 => x"87c9e9fe",
  1898 => x"497086c4",
  1899 => x"eac00299",
  1900 => x"a61ec487",
  1901 => x"f8c21e4d",
  1902 => x"eefe49fc",
  1903 => x"86c887fe",
  1904 => x"d6029870",
  1905 => x"c14a7587",
  1906 => x"c449d1f8",
  1907 => x"d9cafe4b",
  1908 => x"02987087",
  1909 => x"48c087ca",
  1910 => x"c087edc0",
  1911 => x"87e8c048",
  1912 => x"c187f3c0",
  1913 => x"987087c4",
  1914 => x"c087c802",
  1915 => x"987087fc",
  1916 => x"c287f805",
  1917 => x"02bfdcf9",
  1918 => x"f8c287cc",
  1919 => x"f9c248f8",
  1920 => x"fc78bfdc",
  1921 => x"48c187d4",
  1922 => x"264d2626",
  1923 => x"264b264c",
  1924 => x"52415b4f",
  1925 => x"c01e0043",
  1926 => x"fcf8c21e",
  1927 => x"f4ebfe49",
  1928 => x"d4f9c287",
  1929 => x"2678c048",
  1930 => x"5e0e4f26",
  1931 => x"0e5d5c5b",
  1932 => x"a6c486f4",
  1933 => x"c278c048",
  1934 => x"48bfd4f9",
  1935 => x"03a8b7c3",
  1936 => x"f9c287d1",
  1937 => x"c148bfd4",
  1938 => x"d8f9c280",
  1939 => x"48fbc058",
  1940 => x"c287e2c6",
  1941 => x"fe49fcf8",
  1942 => x"7087f5f0",
  1943 => x"d4f9c24c",
  1944 => x"8ac34abf",
  1945 => x"c187d802",
  1946 => x"cbc5028a",
  1947 => x"c2028a87",
  1948 => x"028a87f6",
  1949 => x"8a87cdc1",
  1950 => x"87e2c302",
  1951 => x"c087e1c5",
  1952 => x"c44a754d",
  1953 => x"d3c0c292",
  1954 => x"d0f9c282",
  1955 => x"70807548",
  1956 => x"bf976e7e",
  1957 => x"6e4b494b",
  1958 => x"50a3c148",
  1959 => x"4811816a",
  1960 => x"7058a6cc",
  1961 => x"87c402ac",
  1962 => x"50c0486e",
  1963 => x"c70566c8",
  1964 => x"d4f9c287",
  1965 => x"78a5c448",
  1966 => x"b7c485c1",
  1967 => x"c0ff04ad",
  1968 => x"87dcc487",
  1969 => x"bfe0f9c2",
  1970 => x"a8b7c848",
  1971 => x"ca87d101",
  1972 => x"87cc02ac",
  1973 => x"c702accd",
  1974 => x"acb7c087",
  1975 => x"87f3c003",
  1976 => x"bfe0f9c2",
  1977 => x"abb7c84b",
  1978 => x"c287d203",
  1979 => x"7349e4f9",
  1980 => x"51e0c081",
  1981 => x"b7c883c1",
  1982 => x"eeff04ab",
  1983 => x"ecf9c287",
  1984 => x"50d2c148",
  1985 => x"c150cfc1",
  1986 => x"50c050cd",
  1987 => x"78c380e4",
  1988 => x"c287cdc3",
  1989 => x"49bfe0f9",
  1990 => x"c280c148",
  1991 => x"4858e4f9",
  1992 => x"7481a0c4",
  1993 => x"87f8c251",
  1994 => x"acb7f0c0",
  1995 => x"c087da04",
  1996 => x"01acb7f9",
  1997 => x"f9c287d3",
  1998 => x"ca49bfd8",
  1999 => x"c04a7491",
  2000 => x"f9c28af0",
  2001 => x"a17248d8",
  2002 => x"02acca78",
  2003 => x"cd87c6c0",
  2004 => x"cbc205ac",
  2005 => x"d4f9c287",
  2006 => x"c278c348",
  2007 => x"f0c087c2",
  2008 => x"db04acb7",
  2009 => x"b7f9c087",
  2010 => x"d3c001ac",
  2011 => x"dcf9c287",
  2012 => x"91d049bf",
  2013 => x"f0c04a74",
  2014 => x"dcf9c28a",
  2015 => x"78a17248",
  2016 => x"acb7c1c1",
  2017 => x"87dbc004",
  2018 => x"acb7c6c1",
  2019 => x"87d3c001",
  2020 => x"bfdcf9c2",
  2021 => x"7491d049",
  2022 => x"8af7c04a",
  2023 => x"48dcf9c2",
  2024 => x"ca78a172",
  2025 => x"c6c002ac",
  2026 => x"05accd87",
  2027 => x"c287f1c0",
  2028 => x"c348d4f9",
  2029 => x"87e8c078",
  2030 => x"05ace2c0",
  2031 => x"c487c9c0",
  2032 => x"fbc048a6",
  2033 => x"87d8c078",
  2034 => x"c002acca",
  2035 => x"accd87c6",
  2036 => x"87c9c005",
  2037 => x"48d4f9c2",
  2038 => x"c3c078c3",
  2039 => x"5ca6c887",
  2040 => x"03acb7c0",
  2041 => x"4887c4c0",
  2042 => x"c487cac0",
  2043 => x"c6f90266",
  2044 => x"ffc34887",
  2045 => x"f88ef499",
  2046 => x"4f4387cf",
  2047 => x"003d464e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
