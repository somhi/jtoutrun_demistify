
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"fc",x"f7",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"fc",x"f7",x"c2"),
    14 => (x"48",x"fc",x"e4",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e6",x"e5"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"81",x"48",x"73",x"1e"),
    47 => (x"72",x"05",x"a9",x"73"),
    48 => (x"26",x"87",x"f9",x"53"),
    49 => (x"4a",x"71",x"1e",x"4f"),
    50 => (x"48",x"49",x"66",x"c4"),
    51 => (x"a6",x"c8",x"88",x"c1"),
    52 => (x"02",x"99",x"71",x"58"),
    53 => (x"d4",x"ff",x"87",x"d6"),
    54 => (x"78",x"ff",x"c3",x"48"),
    55 => (x"66",x"c4",x"52",x"68"),
    56 => (x"88",x"c1",x"48",x"49"),
    57 => (x"71",x"58",x"a6",x"c8"),
    58 => (x"87",x"ea",x"05",x"99"),
    59 => (x"73",x"1e",x"4f",x"26"),
    60 => (x"4b",x"d4",x"ff",x"1e"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"7b",x"ff",x"c3",x"4a"),
    63 => (x"32",x"c8",x"49",x"6b"),
    64 => (x"ff",x"c3",x"b1",x"72"),
    65 => (x"c8",x"4a",x"6b",x"7b"),
    66 => (x"c3",x"b2",x"71",x"31"),
    67 => (x"49",x"6b",x"7b",x"ff"),
    68 => (x"b1",x"72",x"32",x"c8"),
    69 => (x"87",x"c4",x"48",x"71"),
    70 => (x"4c",x"26",x"4d",x"26"),
    71 => (x"4f",x"26",x"4b",x"26"),
    72 => (x"5c",x"5b",x"5e",x"0e"),
    73 => (x"4a",x"71",x"0e",x"5d"),
    74 => (x"72",x"4c",x"d4",x"ff"),
    75 => (x"99",x"ff",x"c3",x"49"),
    76 => (x"e4",x"c2",x"7c",x"71"),
    77 => (x"c8",x"05",x"bf",x"fc"),
    78 => (x"48",x"66",x"d0",x"87"),
    79 => (x"a6",x"d4",x"30",x"c9"),
    80 => (x"49",x"66",x"d0",x"58"),
    81 => (x"ff",x"c3",x"29",x"d8"),
    82 => (x"d0",x"7c",x"71",x"99"),
    83 => (x"29",x"d0",x"49",x"66"),
    84 => (x"71",x"99",x"ff",x"c3"),
    85 => (x"49",x"66",x"d0",x"7c"),
    86 => (x"ff",x"c3",x"29",x"c8"),
    87 => (x"d0",x"7c",x"71",x"99"),
    88 => (x"ff",x"c3",x"49",x"66"),
    89 => (x"72",x"7c",x"71",x"99"),
    90 => (x"c3",x"29",x"d0",x"49"),
    91 => (x"7c",x"71",x"99",x"ff"),
    92 => (x"f0",x"c9",x"4b",x"6c"),
    93 => (x"ff",x"c3",x"4d",x"ff"),
    94 => (x"87",x"d0",x"05",x"ab"),
    95 => (x"6c",x"7c",x"ff",x"c3"),
    96 => (x"02",x"8d",x"c1",x"4b"),
    97 => (x"ff",x"c3",x"87",x"c6"),
    98 => (x"87",x"f0",x"02",x"ab"),
    99 => (x"c7",x"fe",x"48",x"73"),
   100 => (x"49",x"c0",x"1e",x"87"),
   101 => (x"c3",x"48",x"d4",x"ff"),
   102 => (x"81",x"c1",x"78",x"ff"),
   103 => (x"a9",x"b7",x"c8",x"c3"),
   104 => (x"26",x"87",x"f1",x"04"),
   105 => (x"1e",x"73",x"1e",x"4f"),
   106 => (x"f8",x"c4",x"87",x"e7"),
   107 => (x"1e",x"c0",x"4b",x"df"),
   108 => (x"c1",x"f0",x"ff",x"c0"),
   109 => (x"e7",x"fd",x"49",x"f7"),
   110 => (x"c1",x"86",x"c4",x"87"),
   111 => (x"ea",x"c0",x"05",x"a8"),
   112 => (x"48",x"d4",x"ff",x"87"),
   113 => (x"c1",x"78",x"ff",x"c3"),
   114 => (x"c0",x"c0",x"c0",x"c0"),
   115 => (x"e1",x"c0",x"1e",x"c0"),
   116 => (x"49",x"e9",x"c1",x"f0"),
   117 => (x"c4",x"87",x"c9",x"fd"),
   118 => (x"05",x"98",x"70",x"86"),
   119 => (x"d4",x"ff",x"87",x"ca"),
   120 => (x"78",x"ff",x"c3",x"48"),
   121 => (x"87",x"cb",x"48",x"c1"),
   122 => (x"c1",x"87",x"e6",x"fe"),
   123 => (x"fd",x"fe",x"05",x"8b"),
   124 => (x"fc",x"48",x"c0",x"87"),
   125 => (x"73",x"1e",x"87",x"e6"),
   126 => (x"48",x"d4",x"ff",x"1e"),
   127 => (x"d3",x"78",x"ff",x"c3"),
   128 => (x"c0",x"1e",x"c0",x"4b"),
   129 => (x"c1",x"c1",x"f0",x"ff"),
   130 => (x"87",x"d4",x"fc",x"49"),
   131 => (x"98",x"70",x"86",x"c4"),
   132 => (x"ff",x"87",x"ca",x"05"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"cb",x"48",x"c1",x"78"),
   135 => (x"87",x"f1",x"fd",x"87"),
   136 => (x"ff",x"05",x"8b",x"c1"),
   137 => (x"48",x"c0",x"87",x"db"),
   138 => (x"0e",x"87",x"f1",x"fb"),
   139 => (x"0e",x"5c",x"5b",x"5e"),
   140 => (x"fd",x"4c",x"d4",x"ff"),
   141 => (x"ea",x"c6",x"87",x"db"),
   142 => (x"f0",x"e1",x"c0",x"1e"),
   143 => (x"fb",x"49",x"c8",x"c1"),
   144 => (x"86",x"c4",x"87",x"de"),
   145 => (x"c8",x"02",x"a8",x"c1"),
   146 => (x"87",x"ea",x"fe",x"87"),
   147 => (x"e2",x"c1",x"48",x"c0"),
   148 => (x"87",x"da",x"fa",x"87"),
   149 => (x"ff",x"cf",x"49",x"70"),
   150 => (x"ea",x"c6",x"99",x"ff"),
   151 => (x"87",x"c8",x"02",x"a9"),
   152 => (x"c0",x"87",x"d3",x"fe"),
   153 => (x"87",x"cb",x"c1",x"48"),
   154 => (x"c0",x"7c",x"ff",x"c3"),
   155 => (x"f4",x"fc",x"4b",x"f1"),
   156 => (x"02",x"98",x"70",x"87"),
   157 => (x"c0",x"87",x"eb",x"c0"),
   158 => (x"f0",x"ff",x"c0",x"1e"),
   159 => (x"fa",x"49",x"fa",x"c1"),
   160 => (x"86",x"c4",x"87",x"de"),
   161 => (x"d9",x"05",x"98",x"70"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"ff",x"c3",x"49",x"6c"),
   164 => (x"7c",x"7c",x"7c",x"7c"),
   165 => (x"02",x"99",x"c0",x"c1"),
   166 => (x"48",x"c1",x"87",x"c4"),
   167 => (x"48",x"c0",x"87",x"d5"),
   168 => (x"ab",x"c2",x"87",x"d1"),
   169 => (x"c0",x"87",x"c4",x"05"),
   170 => (x"c1",x"87",x"c8",x"48"),
   171 => (x"fd",x"fe",x"05",x"8b"),
   172 => (x"f9",x"48",x"c0",x"87"),
   173 => (x"73",x"1e",x"87",x"e4"),
   174 => (x"fc",x"e4",x"c2",x"1e"),
   175 => (x"c7",x"78",x"c1",x"48"),
   176 => (x"48",x"d0",x"ff",x"4b"),
   177 => (x"c8",x"fb",x"78",x"c2"),
   178 => (x"48",x"d0",x"ff",x"87"),
   179 => (x"1e",x"c0",x"78",x"c3"),
   180 => (x"c1",x"d0",x"e5",x"c0"),
   181 => (x"c7",x"f9",x"49",x"c0"),
   182 => (x"c1",x"86",x"c4",x"87"),
   183 => (x"87",x"c1",x"05",x"a8"),
   184 => (x"05",x"ab",x"c2",x"4b"),
   185 => (x"48",x"c0",x"87",x"c5"),
   186 => (x"c1",x"87",x"f9",x"c0"),
   187 => (x"d0",x"ff",x"05",x"8b"),
   188 => (x"87",x"f7",x"fc",x"87"),
   189 => (x"58",x"c0",x"e5",x"c2"),
   190 => (x"cd",x"05",x"98",x"70"),
   191 => (x"c0",x"1e",x"c1",x"87"),
   192 => (x"d0",x"c1",x"f0",x"ff"),
   193 => (x"87",x"d8",x"f8",x"49"),
   194 => (x"d4",x"ff",x"86",x"c4"),
   195 => (x"78",x"ff",x"c3",x"48"),
   196 => (x"c2",x"87",x"fc",x"c2"),
   197 => (x"ff",x"58",x"c4",x"e5"),
   198 => (x"78",x"c2",x"48",x"d0"),
   199 => (x"c3",x"48",x"d4",x"ff"),
   200 => (x"48",x"c1",x"78",x"ff"),
   201 => (x"0e",x"87",x"f5",x"f7"),
   202 => (x"5d",x"5c",x"5b",x"5e"),
   203 => (x"c0",x"4b",x"71",x"0e"),
   204 => (x"cd",x"ee",x"c5",x"4c"),
   205 => (x"d4",x"ff",x"4a",x"df"),
   206 => (x"78",x"ff",x"c3",x"48"),
   207 => (x"fe",x"c3",x"49",x"68"),
   208 => (x"fd",x"c0",x"05",x"a9"),
   209 => (x"73",x"4d",x"70",x"87"),
   210 => (x"87",x"cc",x"02",x"9b"),
   211 => (x"73",x"1e",x"66",x"d0"),
   212 => (x"87",x"f1",x"f5",x"49"),
   213 => (x"87",x"d6",x"86",x"c4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"ff",x"c3",x"78",x"d1"),
   216 => (x"48",x"66",x"d0",x"7d"),
   217 => (x"a6",x"d4",x"88",x"c1"),
   218 => (x"05",x"98",x"70",x"58"),
   219 => (x"d4",x"ff",x"87",x"f0"),
   220 => (x"78",x"ff",x"c3",x"48"),
   221 => (x"05",x"9b",x"73",x"78"),
   222 => (x"d0",x"ff",x"87",x"c5"),
   223 => (x"c1",x"78",x"d0",x"48"),
   224 => (x"8a",x"c1",x"4c",x"4a"),
   225 => (x"87",x"ee",x"fe",x"05"),
   226 => (x"cb",x"f6",x"48",x"74"),
   227 => (x"1e",x"73",x"1e",x"87"),
   228 => (x"4b",x"c0",x"4a",x"71"),
   229 => (x"c3",x"48",x"d4",x"ff"),
   230 => (x"d0",x"ff",x"78",x"ff"),
   231 => (x"78",x"c3",x"c4",x"48"),
   232 => (x"c3",x"48",x"d4",x"ff"),
   233 => (x"1e",x"72",x"78",x"ff"),
   234 => (x"c1",x"f0",x"ff",x"c0"),
   235 => (x"ef",x"f5",x"49",x"d1"),
   236 => (x"70",x"86",x"c4",x"87"),
   237 => (x"87",x"d2",x"05",x"98"),
   238 => (x"cc",x"1e",x"c0",x"c8"),
   239 => (x"e6",x"fd",x"49",x"66"),
   240 => (x"70",x"86",x"c4",x"87"),
   241 => (x"48",x"d0",x"ff",x"4b"),
   242 => (x"48",x"73",x"78",x"c2"),
   243 => (x"0e",x"87",x"cd",x"f5"),
   244 => (x"5d",x"5c",x"5b",x"5e"),
   245 => (x"c0",x"1e",x"c0",x"0e"),
   246 => (x"c9",x"c1",x"f0",x"ff"),
   247 => (x"87",x"c0",x"f5",x"49"),
   248 => (x"e5",x"c2",x"1e",x"d2"),
   249 => (x"fe",x"fc",x"49",x"c4"),
   250 => (x"c0",x"86",x"c8",x"87"),
   251 => (x"d2",x"84",x"c1",x"4c"),
   252 => (x"f8",x"04",x"ac",x"b7"),
   253 => (x"c4",x"e5",x"c2",x"87"),
   254 => (x"c3",x"49",x"bf",x"97"),
   255 => (x"c0",x"c1",x"99",x"c0"),
   256 => (x"e7",x"c0",x"05",x"a9"),
   257 => (x"cb",x"e5",x"c2",x"87"),
   258 => (x"d0",x"49",x"bf",x"97"),
   259 => (x"cc",x"e5",x"c2",x"31"),
   260 => (x"c8",x"4a",x"bf",x"97"),
   261 => (x"c2",x"b1",x"72",x"32"),
   262 => (x"bf",x"97",x"cd",x"e5"),
   263 => (x"4c",x"71",x"b1",x"4a"),
   264 => (x"ff",x"ff",x"ff",x"cf"),
   265 => (x"ca",x"84",x"c1",x"9c"),
   266 => (x"87",x"e7",x"c1",x"34"),
   267 => (x"97",x"cd",x"e5",x"c2"),
   268 => (x"31",x"c1",x"49",x"bf"),
   269 => (x"e5",x"c2",x"99",x"c6"),
   270 => (x"4a",x"bf",x"97",x"ce"),
   271 => (x"72",x"2a",x"b7",x"c7"),
   272 => (x"c9",x"e5",x"c2",x"b1"),
   273 => (x"4d",x"4a",x"bf",x"97"),
   274 => (x"e5",x"c2",x"9d",x"cf"),
   275 => (x"4a",x"bf",x"97",x"ca"),
   276 => (x"32",x"ca",x"9a",x"c3"),
   277 => (x"97",x"cb",x"e5",x"c2"),
   278 => (x"33",x"c2",x"4b",x"bf"),
   279 => (x"e5",x"c2",x"b2",x"73"),
   280 => (x"4b",x"bf",x"97",x"cc"),
   281 => (x"c6",x"9b",x"c0",x"c3"),
   282 => (x"b2",x"73",x"2b",x"b7"),
   283 => (x"48",x"c1",x"81",x"c2"),
   284 => (x"49",x"70",x"30",x"71"),
   285 => (x"30",x"75",x"48",x"c1"),
   286 => (x"4c",x"72",x"4d",x"70"),
   287 => (x"94",x"71",x"84",x"c1"),
   288 => (x"ad",x"b7",x"c0",x"c8"),
   289 => (x"c1",x"87",x"cc",x"06"),
   290 => (x"c8",x"2d",x"b7",x"34"),
   291 => (x"01",x"ad",x"b7",x"c0"),
   292 => (x"74",x"87",x"f4",x"ff"),
   293 => (x"87",x"c0",x"f2",x"48"),
   294 => (x"5c",x"5b",x"5e",x"0e"),
   295 => (x"86",x"f8",x"0e",x"5d"),
   296 => (x"48",x"ea",x"ed",x"c2"),
   297 => (x"e5",x"c2",x"78",x"c0"),
   298 => (x"49",x"c0",x"1e",x"e2"),
   299 => (x"c4",x"87",x"de",x"fb"),
   300 => (x"05",x"98",x"70",x"86"),
   301 => (x"48",x"c0",x"87",x"c5"),
   302 => (x"c0",x"87",x"ce",x"c9"),
   303 => (x"c0",x"7e",x"c1",x"4d"),
   304 => (x"49",x"bf",x"d8",x"f5"),
   305 => (x"4a",x"d8",x"e6",x"c2"),
   306 => (x"ee",x"4b",x"c8",x"71"),
   307 => (x"98",x"70",x"87",x"dc"),
   308 => (x"c0",x"87",x"c2",x"05"),
   309 => (x"d4",x"f5",x"c0",x"7e"),
   310 => (x"e6",x"c2",x"49",x"bf"),
   311 => (x"c8",x"71",x"4a",x"f4"),
   312 => (x"87",x"c6",x"ee",x"4b"),
   313 => (x"c2",x"05",x"98",x"70"),
   314 => (x"6e",x"7e",x"c0",x"87"),
   315 => (x"87",x"fd",x"c0",x"02"),
   316 => (x"bf",x"e8",x"ec",x"c2"),
   317 => (x"e0",x"ed",x"c2",x"4d"),
   318 => (x"48",x"7e",x"bf",x"9f"),
   319 => (x"a8",x"ea",x"d6",x"c5"),
   320 => (x"c2",x"87",x"c7",x"05"),
   321 => (x"4d",x"bf",x"e8",x"ec"),
   322 => (x"48",x"6e",x"87",x"ce"),
   323 => (x"a8",x"d5",x"e9",x"ca"),
   324 => (x"c0",x"87",x"c5",x"02"),
   325 => (x"87",x"f1",x"c7",x"48"),
   326 => (x"1e",x"e2",x"e5",x"c2"),
   327 => (x"ec",x"f9",x"49",x"75"),
   328 => (x"70",x"86",x"c4",x"87"),
   329 => (x"87",x"c5",x"05",x"98"),
   330 => (x"dc",x"c7",x"48",x"c0"),
   331 => (x"d4",x"f5",x"c0",x"87"),
   332 => (x"e6",x"c2",x"49",x"bf"),
   333 => (x"c8",x"71",x"4a",x"f4"),
   334 => (x"87",x"ee",x"ec",x"4b"),
   335 => (x"c8",x"05",x"98",x"70"),
   336 => (x"ea",x"ed",x"c2",x"87"),
   337 => (x"da",x"78",x"c1",x"48"),
   338 => (x"d8",x"f5",x"c0",x"87"),
   339 => (x"e6",x"c2",x"49",x"bf"),
   340 => (x"c8",x"71",x"4a",x"d8"),
   341 => (x"87",x"d2",x"ec",x"4b"),
   342 => (x"c0",x"02",x"98",x"70"),
   343 => (x"48",x"c0",x"87",x"c5"),
   344 => (x"c2",x"87",x"e6",x"c6"),
   345 => (x"bf",x"97",x"e0",x"ed"),
   346 => (x"a9",x"d5",x"c1",x"49"),
   347 => (x"87",x"cd",x"c0",x"05"),
   348 => (x"97",x"e1",x"ed",x"c2"),
   349 => (x"ea",x"c2",x"49",x"bf"),
   350 => (x"c5",x"c0",x"02",x"a9"),
   351 => (x"c6",x"48",x"c0",x"87"),
   352 => (x"e5",x"c2",x"87",x"c7"),
   353 => (x"7e",x"bf",x"97",x"e2"),
   354 => (x"a8",x"e9",x"c3",x"48"),
   355 => (x"87",x"ce",x"c0",x"02"),
   356 => (x"eb",x"c3",x"48",x"6e"),
   357 => (x"c5",x"c0",x"02",x"a8"),
   358 => (x"c5",x"48",x"c0",x"87"),
   359 => (x"e5",x"c2",x"87",x"eb"),
   360 => (x"49",x"bf",x"97",x"ed"),
   361 => (x"cc",x"c0",x"05",x"99"),
   362 => (x"ee",x"e5",x"c2",x"87"),
   363 => (x"c2",x"49",x"bf",x"97"),
   364 => (x"c5",x"c0",x"02",x"a9"),
   365 => (x"c5",x"48",x"c0",x"87"),
   366 => (x"e5",x"c2",x"87",x"cf"),
   367 => (x"48",x"bf",x"97",x"ef"),
   368 => (x"58",x"e6",x"ed",x"c2"),
   369 => (x"c1",x"48",x"4c",x"70"),
   370 => (x"ea",x"ed",x"c2",x"88"),
   371 => (x"f0",x"e5",x"c2",x"58"),
   372 => (x"75",x"49",x"bf",x"97"),
   373 => (x"f1",x"e5",x"c2",x"81"),
   374 => (x"c8",x"4a",x"bf",x"97"),
   375 => (x"7e",x"a1",x"72",x"32"),
   376 => (x"48",x"f7",x"f1",x"c2"),
   377 => (x"e5",x"c2",x"78",x"6e"),
   378 => (x"48",x"bf",x"97",x"f2"),
   379 => (x"c2",x"58",x"a6",x"c8"),
   380 => (x"02",x"bf",x"ea",x"ed"),
   381 => (x"c0",x"87",x"d4",x"c2"),
   382 => (x"49",x"bf",x"d4",x"f5"),
   383 => (x"4a",x"f4",x"e6",x"c2"),
   384 => (x"e9",x"4b",x"c8",x"71"),
   385 => (x"98",x"70",x"87",x"e4"),
   386 => (x"87",x"c5",x"c0",x"02"),
   387 => (x"f8",x"c3",x"48",x"c0"),
   388 => (x"e2",x"ed",x"c2",x"87"),
   389 => (x"f2",x"c2",x"4c",x"bf"),
   390 => (x"e6",x"c2",x"5c",x"cb"),
   391 => (x"49",x"bf",x"97",x"c7"),
   392 => (x"e6",x"c2",x"31",x"c8"),
   393 => (x"4a",x"bf",x"97",x"c6"),
   394 => (x"e6",x"c2",x"49",x"a1"),
   395 => (x"4a",x"bf",x"97",x"c8"),
   396 => (x"a1",x"72",x"32",x"d0"),
   397 => (x"c9",x"e6",x"c2",x"49"),
   398 => (x"d8",x"4a",x"bf",x"97"),
   399 => (x"49",x"a1",x"72",x"32"),
   400 => (x"c2",x"91",x"66",x"c4"),
   401 => (x"81",x"bf",x"f7",x"f1"),
   402 => (x"59",x"ff",x"f1",x"c2"),
   403 => (x"97",x"cf",x"e6",x"c2"),
   404 => (x"32",x"c8",x"4a",x"bf"),
   405 => (x"97",x"ce",x"e6",x"c2"),
   406 => (x"4a",x"a2",x"4b",x"bf"),
   407 => (x"97",x"d0",x"e6",x"c2"),
   408 => (x"33",x"d0",x"4b",x"bf"),
   409 => (x"c2",x"4a",x"a2",x"73"),
   410 => (x"bf",x"97",x"d1",x"e6"),
   411 => (x"d8",x"9b",x"cf",x"4b"),
   412 => (x"4a",x"a2",x"73",x"33"),
   413 => (x"5a",x"c3",x"f2",x"c2"),
   414 => (x"bf",x"ff",x"f1",x"c2"),
   415 => (x"74",x"8a",x"c2",x"4a"),
   416 => (x"c3",x"f2",x"c2",x"92"),
   417 => (x"78",x"a1",x"72",x"48"),
   418 => (x"c2",x"87",x"ca",x"c1"),
   419 => (x"bf",x"97",x"f4",x"e5"),
   420 => (x"c2",x"31",x"c8",x"49"),
   421 => (x"bf",x"97",x"f3",x"e5"),
   422 => (x"c2",x"49",x"a1",x"4a"),
   423 => (x"c2",x"59",x"f2",x"ed"),
   424 => (x"49",x"bf",x"ee",x"ed"),
   425 => (x"ff",x"c7",x"31",x"c5"),
   426 => (x"c2",x"29",x"c9",x"81"),
   427 => (x"c2",x"59",x"cb",x"f2"),
   428 => (x"bf",x"97",x"f9",x"e5"),
   429 => (x"c2",x"32",x"c8",x"4a"),
   430 => (x"bf",x"97",x"f8",x"e5"),
   431 => (x"c4",x"4a",x"a2",x"4b"),
   432 => (x"82",x"6e",x"92",x"66"),
   433 => (x"5a",x"c7",x"f2",x"c2"),
   434 => (x"48",x"ff",x"f1",x"c2"),
   435 => (x"f1",x"c2",x"78",x"c0"),
   436 => (x"a1",x"72",x"48",x"fb"),
   437 => (x"cb",x"f2",x"c2",x"78"),
   438 => (x"ff",x"f1",x"c2",x"48"),
   439 => (x"f2",x"c2",x"78",x"bf"),
   440 => (x"f2",x"c2",x"48",x"cf"),
   441 => (x"c2",x"78",x"bf",x"c3"),
   442 => (x"02",x"bf",x"ea",x"ed"),
   443 => (x"74",x"87",x"c9",x"c0"),
   444 => (x"70",x"30",x"c4",x"48"),
   445 => (x"87",x"c9",x"c0",x"7e"),
   446 => (x"bf",x"c7",x"f2",x"c2"),
   447 => (x"70",x"30",x"c4",x"48"),
   448 => (x"ee",x"ed",x"c2",x"7e"),
   449 => (x"c1",x"78",x"6e",x"48"),
   450 => (x"26",x"8e",x"f8",x"48"),
   451 => (x"26",x"4c",x"26",x"4d"),
   452 => (x"0e",x"4f",x"26",x"4b"),
   453 => (x"5d",x"5c",x"5b",x"5e"),
   454 => (x"c2",x"4a",x"71",x"0e"),
   455 => (x"02",x"bf",x"ea",x"ed"),
   456 => (x"4b",x"72",x"87",x"cb"),
   457 => (x"4c",x"72",x"2b",x"c7"),
   458 => (x"c9",x"9c",x"ff",x"c1"),
   459 => (x"c8",x"4b",x"72",x"87"),
   460 => (x"c3",x"4c",x"72",x"2b"),
   461 => (x"f1",x"c2",x"9c",x"ff"),
   462 => (x"c0",x"83",x"bf",x"f7"),
   463 => (x"ab",x"bf",x"d0",x"f5"),
   464 => (x"c0",x"87",x"d9",x"02"),
   465 => (x"c2",x"5b",x"d4",x"f5"),
   466 => (x"73",x"1e",x"e2",x"e5"),
   467 => (x"87",x"fd",x"f0",x"49"),
   468 => (x"98",x"70",x"86",x"c4"),
   469 => (x"c0",x"87",x"c5",x"05"),
   470 => (x"87",x"e6",x"c0",x"48"),
   471 => (x"bf",x"ea",x"ed",x"c2"),
   472 => (x"74",x"87",x"d2",x"02"),
   473 => (x"c2",x"91",x"c4",x"49"),
   474 => (x"69",x"81",x"e2",x"e5"),
   475 => (x"ff",x"ff",x"cf",x"4d"),
   476 => (x"cb",x"9d",x"ff",x"ff"),
   477 => (x"c2",x"49",x"74",x"87"),
   478 => (x"e2",x"e5",x"c2",x"91"),
   479 => (x"4d",x"69",x"9f",x"81"),
   480 => (x"c6",x"fe",x"48",x"75"),
   481 => (x"5b",x"5e",x"0e",x"87"),
   482 => (x"f8",x"0e",x"5d",x"5c"),
   483 => (x"9c",x"4c",x"71",x"86"),
   484 => (x"c0",x"87",x"c5",x"05"),
   485 => (x"87",x"c1",x"c3",x"48"),
   486 => (x"6e",x"7e",x"a4",x"c8"),
   487 => (x"d8",x"78",x"c0",x"48"),
   488 => (x"87",x"c7",x"02",x"66"),
   489 => (x"bf",x"97",x"66",x"d8"),
   490 => (x"c0",x"87",x"c5",x"05"),
   491 => (x"87",x"e9",x"c2",x"48"),
   492 => (x"49",x"c1",x"1e",x"c0"),
   493 => (x"c4",x"87",x"fd",x"ce"),
   494 => (x"9d",x"4d",x"70",x"86"),
   495 => (x"87",x"c2",x"c1",x"02"),
   496 => (x"4a",x"f2",x"ed",x"c2"),
   497 => (x"e2",x"49",x"66",x"d8"),
   498 => (x"98",x"70",x"87",x"c5"),
   499 => (x"87",x"f2",x"c0",x"02"),
   500 => (x"66",x"d8",x"4a",x"75"),
   501 => (x"e2",x"4b",x"cb",x"49"),
   502 => (x"98",x"70",x"87",x"ea"),
   503 => (x"87",x"e2",x"c0",x"02"),
   504 => (x"9d",x"75",x"1e",x"c0"),
   505 => (x"c8",x"87",x"c7",x"02"),
   506 => (x"78",x"c0",x"48",x"a6"),
   507 => (x"a6",x"c8",x"87",x"c5"),
   508 => (x"c8",x"78",x"c1",x"48"),
   509 => (x"fb",x"cd",x"49",x"66"),
   510 => (x"70",x"86",x"c4",x"87"),
   511 => (x"fe",x"05",x"9d",x"4d"),
   512 => (x"9d",x"75",x"87",x"fe"),
   513 => (x"87",x"cf",x"c1",x"02"),
   514 => (x"6e",x"49",x"a5",x"dc"),
   515 => (x"da",x"78",x"69",x"48"),
   516 => (x"a6",x"c4",x"49",x"a5"),
   517 => (x"78",x"a4",x"c4",x"48"),
   518 => (x"c4",x"48",x"69",x"9f"),
   519 => (x"c2",x"78",x"08",x"66"),
   520 => (x"02",x"bf",x"ea",x"ed"),
   521 => (x"a5",x"d4",x"87",x"d2"),
   522 => (x"49",x"69",x"9f",x"49"),
   523 => (x"99",x"ff",x"ff",x"c0"),
   524 => (x"30",x"d0",x"48",x"71"),
   525 => (x"87",x"c2",x"7e",x"70"),
   526 => (x"49",x"6e",x"7e",x"c0"),
   527 => (x"bf",x"66",x"c4",x"48"),
   528 => (x"08",x"66",x"c4",x"80"),
   529 => (x"cc",x"7c",x"c0",x"78"),
   530 => (x"66",x"c4",x"49",x"a4"),
   531 => (x"a4",x"d0",x"79",x"bf"),
   532 => (x"c1",x"79",x"c0",x"49"),
   533 => (x"c0",x"87",x"c2",x"48"),
   534 => (x"fa",x"8e",x"f8",x"48"),
   535 => (x"5e",x"0e",x"87",x"ed"),
   536 => (x"0e",x"5d",x"5c",x"5b"),
   537 => (x"02",x"9c",x"4c",x"71"),
   538 => (x"c8",x"87",x"ca",x"c1"),
   539 => (x"02",x"69",x"49",x"a4"),
   540 => (x"d0",x"87",x"c2",x"c1"),
   541 => (x"49",x"6c",x"4a",x"66"),
   542 => (x"5a",x"a6",x"d4",x"82"),
   543 => (x"b9",x"4d",x"66",x"d0"),
   544 => (x"bf",x"e6",x"ed",x"c2"),
   545 => (x"72",x"ba",x"ff",x"4a"),
   546 => (x"02",x"99",x"71",x"99"),
   547 => (x"c4",x"87",x"e4",x"c0"),
   548 => (x"49",x"6b",x"4b",x"a4"),
   549 => (x"70",x"87",x"fc",x"f9"),
   550 => (x"e2",x"ed",x"c2",x"7b"),
   551 => (x"81",x"6c",x"49",x"bf"),
   552 => (x"b9",x"75",x"7c",x"71"),
   553 => (x"bf",x"e6",x"ed",x"c2"),
   554 => (x"72",x"ba",x"ff",x"4a"),
   555 => (x"05",x"99",x"71",x"99"),
   556 => (x"75",x"87",x"dc",x"ff"),
   557 => (x"87",x"d3",x"f9",x"7c"),
   558 => (x"71",x"1e",x"73",x"1e"),
   559 => (x"c7",x"02",x"9b",x"4b"),
   560 => (x"49",x"a3",x"c8",x"87"),
   561 => (x"87",x"c5",x"05",x"69"),
   562 => (x"f7",x"c0",x"48",x"c0"),
   563 => (x"fb",x"f1",x"c2",x"87"),
   564 => (x"a3",x"c4",x"4a",x"bf"),
   565 => (x"c2",x"49",x"69",x"49"),
   566 => (x"e2",x"ed",x"c2",x"89"),
   567 => (x"a2",x"71",x"91",x"bf"),
   568 => (x"e6",x"ed",x"c2",x"4a"),
   569 => (x"99",x"6b",x"49",x"bf"),
   570 => (x"c0",x"4a",x"a2",x"71"),
   571 => (x"c8",x"5a",x"d4",x"f5"),
   572 => (x"49",x"72",x"1e",x"66"),
   573 => (x"c4",x"87",x"d6",x"ea"),
   574 => (x"05",x"98",x"70",x"86"),
   575 => (x"48",x"c0",x"87",x"c4"),
   576 => (x"48",x"c1",x"87",x"c2"),
   577 => (x"0e",x"87",x"c8",x"f8"),
   578 => (x"0e",x"5c",x"5b",x"5e"),
   579 => (x"d0",x"4b",x"71",x"1e"),
   580 => (x"2c",x"c9",x"4c",x"66"),
   581 => (x"c1",x"02",x"9b",x"73"),
   582 => (x"a3",x"c8",x"87",x"d4"),
   583 => (x"c1",x"02",x"69",x"49"),
   584 => (x"ed",x"c2",x"87",x"cc"),
   585 => (x"ff",x"49",x"bf",x"e6"),
   586 => (x"99",x"4a",x"6b",x"b9"),
   587 => (x"03",x"ac",x"71",x"7e"),
   588 => (x"7b",x"c0",x"87",x"d1"),
   589 => (x"c0",x"49",x"a3",x"d0"),
   590 => (x"4a",x"a3",x"cc",x"79"),
   591 => (x"6a",x"49",x"a3",x"c4"),
   592 => (x"72",x"87",x"c2",x"79"),
   593 => (x"02",x"9c",x"74",x"8c"),
   594 => (x"49",x"87",x"e3",x"c0"),
   595 => (x"fc",x"49",x"73",x"1e"),
   596 => (x"86",x"c4",x"87",x"cc"),
   597 => (x"c7",x"49",x"66",x"d0"),
   598 => (x"cb",x"02",x"99",x"ff"),
   599 => (x"e2",x"e5",x"c2",x"87"),
   600 => (x"fd",x"49",x"73",x"1e"),
   601 => (x"86",x"c4",x"87",x"d2"),
   602 => (x"d0",x"49",x"a3",x"d0"),
   603 => (x"f6",x"26",x"79",x"66"),
   604 => (x"5e",x"0e",x"87",x"db"),
   605 => (x"0e",x"5d",x"5c",x"5b"),
   606 => (x"a6",x"d0",x"86",x"f0"),
   607 => (x"66",x"e4",x"c0",x"59"),
   608 => (x"02",x"66",x"cc",x"4b"),
   609 => (x"c8",x"48",x"87",x"ca"),
   610 => (x"6e",x"7e",x"70",x"80"),
   611 => (x"87",x"c5",x"05",x"bf"),
   612 => (x"ec",x"c3",x"48",x"c0"),
   613 => (x"4c",x"66",x"cc",x"87"),
   614 => (x"49",x"73",x"84",x"d0"),
   615 => (x"6c",x"48",x"a6",x"c4"),
   616 => (x"81",x"66",x"c4",x"78"),
   617 => (x"bf",x"6e",x"80",x"c4"),
   618 => (x"a9",x"66",x"c8",x"78"),
   619 => (x"49",x"87",x"c6",x"06"),
   620 => (x"71",x"89",x"66",x"c4"),
   621 => (x"ab",x"b7",x"c0",x"4b"),
   622 => (x"48",x"87",x"c4",x"01"),
   623 => (x"c4",x"87",x"c2",x"c3"),
   624 => (x"ff",x"c7",x"48",x"66"),
   625 => (x"6e",x"7e",x"70",x"98"),
   626 => (x"87",x"c9",x"c1",x"02"),
   627 => (x"6e",x"49",x"c0",x"c8"),
   628 => (x"c2",x"4a",x"71",x"89"),
   629 => (x"6e",x"4d",x"e2",x"e5"),
   630 => (x"aa",x"b7",x"73",x"85"),
   631 => (x"4a",x"87",x"c1",x"06"),
   632 => (x"c4",x"48",x"49",x"72"),
   633 => (x"7c",x"70",x"80",x"66"),
   634 => (x"c1",x"49",x"8b",x"72"),
   635 => (x"02",x"99",x"71",x"8a"),
   636 => (x"e0",x"c0",x"87",x"d9"),
   637 => (x"50",x"15",x"48",x"66"),
   638 => (x"48",x"66",x"e0",x"c0"),
   639 => (x"e4",x"c0",x"80",x"c1"),
   640 => (x"49",x"72",x"58",x"a6"),
   641 => (x"99",x"71",x"8a",x"c1"),
   642 => (x"c1",x"87",x"e7",x"05"),
   643 => (x"49",x"66",x"d0",x"1e"),
   644 => (x"c4",x"87",x"cb",x"f9"),
   645 => (x"ab",x"b7",x"c0",x"86"),
   646 => (x"87",x"e3",x"c1",x"06"),
   647 => (x"4d",x"66",x"e0",x"c0"),
   648 => (x"ab",x"b7",x"ff",x"c7"),
   649 => (x"87",x"e2",x"c0",x"06"),
   650 => (x"66",x"d0",x"1e",x"75"),
   651 => (x"87",x"c8",x"fa",x"49"),
   652 => (x"6c",x"85",x"c0",x"c8"),
   653 => (x"80",x"c0",x"c8",x"48"),
   654 => (x"c0",x"c8",x"7c",x"70"),
   655 => (x"d4",x"1e",x"c1",x"8b"),
   656 => (x"d9",x"f8",x"49",x"66"),
   657 => (x"c0",x"86",x"c8",x"87"),
   658 => (x"e5",x"c2",x"87",x"ee"),
   659 => (x"66",x"d0",x"1e",x"e2"),
   660 => (x"87",x"e4",x"f9",x"49"),
   661 => (x"e5",x"c2",x"86",x"c4"),
   662 => (x"49",x"73",x"4a",x"e2"),
   663 => (x"70",x"80",x"6c",x"48"),
   664 => (x"c1",x"49",x"73",x"7c"),
   665 => (x"02",x"99",x"71",x"8b"),
   666 => (x"97",x"12",x"87",x"ce"),
   667 => (x"73",x"85",x"c1",x"7d"),
   668 => (x"71",x"8b",x"c1",x"49"),
   669 => (x"87",x"f2",x"05",x"99"),
   670 => (x"01",x"ab",x"b7",x"c0"),
   671 => (x"c1",x"87",x"e1",x"fe"),
   672 => (x"f2",x"8e",x"f0",x"48"),
   673 => (x"5e",x"0e",x"87",x"c5"),
   674 => (x"0e",x"5d",x"5c",x"5b"),
   675 => (x"02",x"9b",x"4b",x"71"),
   676 => (x"a3",x"c8",x"87",x"c7"),
   677 => (x"c5",x"05",x"6d",x"4d"),
   678 => (x"c0",x"48",x"ff",x"87"),
   679 => (x"a3",x"d0",x"87",x"fd"),
   680 => (x"c7",x"49",x"6c",x"4c"),
   681 => (x"d8",x"05",x"99",x"ff"),
   682 => (x"c9",x"02",x"6c",x"87"),
   683 => (x"73",x"1e",x"c1",x"87"),
   684 => (x"87",x"ea",x"f6",x"49"),
   685 => (x"e5",x"c2",x"86",x"c4"),
   686 => (x"49",x"73",x"1e",x"e2"),
   687 => (x"c4",x"87",x"f9",x"f7"),
   688 => (x"6d",x"4a",x"6c",x"86"),
   689 => (x"87",x"c4",x"04",x"aa"),
   690 => (x"87",x"cf",x"48",x"ff"),
   691 => (x"72",x"7c",x"a2",x"c1"),
   692 => (x"99",x"ff",x"c7",x"49"),
   693 => (x"81",x"e2",x"e5",x"c2"),
   694 => (x"f0",x"48",x"69",x"97"),
   695 => (x"73",x"1e",x"87",x"ed"),
   696 => (x"9b",x"4b",x"71",x"1e"),
   697 => (x"87",x"e4",x"c0",x"02"),
   698 => (x"5b",x"cf",x"f2",x"c2"),
   699 => (x"8a",x"c2",x"4a",x"73"),
   700 => (x"bf",x"e2",x"ed",x"c2"),
   701 => (x"f1",x"c2",x"92",x"49"),
   702 => (x"72",x"48",x"bf",x"fb"),
   703 => (x"d3",x"f2",x"c2",x"80"),
   704 => (x"c4",x"48",x"71",x"58"),
   705 => (x"f2",x"ed",x"c2",x"30"),
   706 => (x"87",x"ed",x"c0",x"58"),
   707 => (x"48",x"cb",x"f2",x"c2"),
   708 => (x"bf",x"ff",x"f1",x"c2"),
   709 => (x"cf",x"f2",x"c2",x"78"),
   710 => (x"c3",x"f2",x"c2",x"48"),
   711 => (x"ed",x"c2",x"78",x"bf"),
   712 => (x"c9",x"02",x"bf",x"ea"),
   713 => (x"e2",x"ed",x"c2",x"87"),
   714 => (x"31",x"c4",x"49",x"bf"),
   715 => (x"f2",x"c2",x"87",x"c7"),
   716 => (x"c4",x"49",x"bf",x"c7"),
   717 => (x"f2",x"ed",x"c2",x"31"),
   718 => (x"87",x"d3",x"ef",x"59"),
   719 => (x"5c",x"5b",x"5e",x"0e"),
   720 => (x"c0",x"4a",x"71",x"0e"),
   721 => (x"02",x"9a",x"72",x"4b"),
   722 => (x"da",x"87",x"e1",x"c0"),
   723 => (x"69",x"9f",x"49",x"a2"),
   724 => (x"ea",x"ed",x"c2",x"4b"),
   725 => (x"87",x"cf",x"02",x"bf"),
   726 => (x"9f",x"49",x"a2",x"d4"),
   727 => (x"c0",x"4c",x"49",x"69"),
   728 => (x"d0",x"9c",x"ff",x"ff"),
   729 => (x"c0",x"87",x"c2",x"34"),
   730 => (x"b3",x"49",x"74",x"4c"),
   731 => (x"ed",x"fd",x"49",x"73"),
   732 => (x"87",x"d9",x"ee",x"87"),
   733 => (x"5c",x"5b",x"5e",x"0e"),
   734 => (x"86",x"f4",x"0e",x"5d"),
   735 => (x"7e",x"c0",x"4a",x"71"),
   736 => (x"d8",x"02",x"9a",x"72"),
   737 => (x"de",x"e5",x"c2",x"87"),
   738 => (x"c2",x"78",x"c0",x"48"),
   739 => (x"c2",x"48",x"d6",x"e5"),
   740 => (x"78",x"bf",x"cf",x"f2"),
   741 => (x"48",x"da",x"e5",x"c2"),
   742 => (x"bf",x"cb",x"f2",x"c2"),
   743 => (x"ff",x"ed",x"c2",x"78"),
   744 => (x"c2",x"50",x"c0",x"48"),
   745 => (x"49",x"bf",x"ee",x"ed"),
   746 => (x"bf",x"de",x"e5",x"c2"),
   747 => (x"03",x"aa",x"71",x"4a"),
   748 => (x"72",x"87",x"ca",x"c4"),
   749 => (x"05",x"99",x"cf",x"49"),
   750 => (x"c0",x"87",x"ea",x"c0"),
   751 => (x"c2",x"48",x"d0",x"f5"),
   752 => (x"78",x"bf",x"d6",x"e5"),
   753 => (x"1e",x"e2",x"e5",x"c2"),
   754 => (x"bf",x"d6",x"e5",x"c2"),
   755 => (x"d6",x"e5",x"c2",x"49"),
   756 => (x"78",x"a1",x"c1",x"48"),
   757 => (x"f4",x"de",x"ff",x"71"),
   758 => (x"c0",x"86",x"c4",x"87"),
   759 => (x"c2",x"48",x"cc",x"f5"),
   760 => (x"cc",x"78",x"e2",x"e5"),
   761 => (x"cc",x"f5",x"c0",x"87"),
   762 => (x"e0",x"c0",x"48",x"bf"),
   763 => (x"d0",x"f5",x"c0",x"80"),
   764 => (x"de",x"e5",x"c2",x"58"),
   765 => (x"80",x"c1",x"48",x"bf"),
   766 => (x"58",x"e2",x"e5",x"c2"),
   767 => (x"00",x"0d",x"4c",x"27"),
   768 => (x"bf",x"97",x"bf",x"00"),
   769 => (x"c2",x"02",x"9d",x"4d"),
   770 => (x"e5",x"c3",x"87",x"e3"),
   771 => (x"dc",x"c2",x"02",x"ad"),
   772 => (x"cc",x"f5",x"c0",x"87"),
   773 => (x"a3",x"cb",x"4b",x"bf"),
   774 => (x"cf",x"4c",x"11",x"49"),
   775 => (x"d2",x"c1",x"05",x"ac"),
   776 => (x"df",x"49",x"75",x"87"),
   777 => (x"cd",x"89",x"c1",x"99"),
   778 => (x"f2",x"ed",x"c2",x"91"),
   779 => (x"4a",x"a3",x"c1",x"81"),
   780 => (x"a3",x"c3",x"51",x"12"),
   781 => (x"c5",x"51",x"12",x"4a"),
   782 => (x"51",x"12",x"4a",x"a3"),
   783 => (x"12",x"4a",x"a3",x"c7"),
   784 => (x"4a",x"a3",x"c9",x"51"),
   785 => (x"a3",x"ce",x"51",x"12"),
   786 => (x"d0",x"51",x"12",x"4a"),
   787 => (x"51",x"12",x"4a",x"a3"),
   788 => (x"12",x"4a",x"a3",x"d2"),
   789 => (x"4a",x"a3",x"d4",x"51"),
   790 => (x"a3",x"d6",x"51",x"12"),
   791 => (x"d8",x"51",x"12",x"4a"),
   792 => (x"51",x"12",x"4a",x"a3"),
   793 => (x"12",x"4a",x"a3",x"dc"),
   794 => (x"4a",x"a3",x"de",x"51"),
   795 => (x"7e",x"c1",x"51",x"12"),
   796 => (x"74",x"87",x"fa",x"c0"),
   797 => (x"05",x"99",x"c8",x"49"),
   798 => (x"74",x"87",x"eb",x"c0"),
   799 => (x"05",x"99",x"d0",x"49"),
   800 => (x"66",x"dc",x"87",x"d1"),
   801 => (x"87",x"cb",x"c0",x"02"),
   802 => (x"66",x"dc",x"49",x"73"),
   803 => (x"02",x"98",x"70",x"0f"),
   804 => (x"6e",x"87",x"d3",x"c0"),
   805 => (x"87",x"c6",x"c0",x"05"),
   806 => (x"48",x"f2",x"ed",x"c2"),
   807 => (x"f5",x"c0",x"50",x"c0"),
   808 => (x"c2",x"48",x"bf",x"cc"),
   809 => (x"ed",x"c2",x"87",x"e1"),
   810 => (x"50",x"c0",x"48",x"ff"),
   811 => (x"ee",x"ed",x"c2",x"7e"),
   812 => (x"e5",x"c2",x"49",x"bf"),
   813 => (x"71",x"4a",x"bf",x"de"),
   814 => (x"f6",x"fb",x"04",x"aa"),
   815 => (x"cf",x"f2",x"c2",x"87"),
   816 => (x"c8",x"c0",x"05",x"bf"),
   817 => (x"ea",x"ed",x"c2",x"87"),
   818 => (x"f8",x"c1",x"02",x"bf"),
   819 => (x"da",x"e5",x"c2",x"87"),
   820 => (x"fe",x"e8",x"49",x"bf"),
   821 => (x"c2",x"49",x"70",x"87"),
   822 => (x"c4",x"59",x"de",x"e5"),
   823 => (x"e5",x"c2",x"48",x"a6"),
   824 => (x"c2",x"78",x"bf",x"da"),
   825 => (x"02",x"bf",x"ea",x"ed"),
   826 => (x"c4",x"87",x"d8",x"c0"),
   827 => (x"ff",x"cf",x"49",x"66"),
   828 => (x"99",x"f8",x"ff",x"ff"),
   829 => (x"c5",x"c0",x"02",x"a9"),
   830 => (x"c0",x"4c",x"c0",x"87"),
   831 => (x"4c",x"c1",x"87",x"e1"),
   832 => (x"c4",x"87",x"dc",x"c0"),
   833 => (x"ff",x"cf",x"49",x"66"),
   834 => (x"02",x"a9",x"99",x"f8"),
   835 => (x"c8",x"87",x"c8",x"c0"),
   836 => (x"78",x"c0",x"48",x"a6"),
   837 => (x"c8",x"87",x"c5",x"c0"),
   838 => (x"78",x"c1",x"48",x"a6"),
   839 => (x"74",x"4c",x"66",x"c8"),
   840 => (x"e0",x"c0",x"05",x"9c"),
   841 => (x"49",x"66",x"c4",x"87"),
   842 => (x"ed",x"c2",x"89",x"c2"),
   843 => (x"91",x"4a",x"bf",x"e2"),
   844 => (x"bf",x"fb",x"f1",x"c2"),
   845 => (x"d6",x"e5",x"c2",x"4a"),
   846 => (x"78",x"a1",x"72",x"48"),
   847 => (x"48",x"de",x"e5",x"c2"),
   848 => (x"de",x"f9",x"78",x"c0"),
   849 => (x"f4",x"48",x"c0",x"87"),
   850 => (x"87",x"ff",x"e6",x"8e"),
   851 => (x"00",x"00",x"00",x"00"),
   852 => (x"ff",x"ff",x"ff",x"ff"),
   853 => (x"00",x"00",x"0d",x"5c"),
   854 => (x"00",x"00",x"0d",x"65"),
   855 => (x"33",x"54",x"41",x"46"),
   856 => (x"20",x"20",x"20",x"32"),
   857 => (x"54",x"41",x"46",x"00"),
   858 => (x"20",x"20",x"36",x"31"),
   859 => (x"c2",x"1e",x"00",x"20"),
   860 => (x"48",x"bf",x"d4",x"f2"),
   861 => (x"c9",x"05",x"a8",x"dd"),
   862 => (x"da",x"c2",x"c1",x"87"),
   863 => (x"4a",x"49",x"70",x"87"),
   864 => (x"d4",x"ff",x"87",x"c8"),
   865 => (x"78",x"ff",x"c3",x"48"),
   866 => (x"48",x"72",x"4a",x"68"),
   867 => (x"c2",x"1e",x"4f",x"26"),
   868 => (x"48",x"bf",x"d4",x"f2"),
   869 => (x"c6",x"05",x"a8",x"dd"),
   870 => (x"e6",x"c1",x"c1",x"87"),
   871 => (x"ff",x"87",x"d9",x"87"),
   872 => (x"ff",x"c3",x"48",x"d4"),
   873 => (x"48",x"d0",x"ff",x"78"),
   874 => (x"ff",x"78",x"e1",x"c0"),
   875 => (x"78",x"d4",x"48",x"d4"),
   876 => (x"48",x"d3",x"f2",x"c2"),
   877 => (x"50",x"bf",x"d4",x"ff"),
   878 => (x"ff",x"1e",x"4f",x"26"),
   879 => (x"e0",x"c0",x"48",x"d0"),
   880 => (x"1e",x"4f",x"26",x"78"),
   881 => (x"70",x"87",x"e7",x"fe"),
   882 => (x"c6",x"02",x"99",x"49"),
   883 => (x"a9",x"fb",x"c0",x"87"),
   884 => (x"71",x"87",x"f1",x"05"),
   885 => (x"0e",x"4f",x"26",x"48"),
   886 => (x"0e",x"5c",x"5b",x"5e"),
   887 => (x"4c",x"c0",x"4b",x"71"),
   888 => (x"70",x"87",x"cb",x"fe"),
   889 => (x"c0",x"02",x"99",x"49"),
   890 => (x"ec",x"c0",x"87",x"f9"),
   891 => (x"f2",x"c0",x"02",x"a9"),
   892 => (x"a9",x"fb",x"c0",x"87"),
   893 => (x"87",x"eb",x"c0",x"02"),
   894 => (x"ac",x"b7",x"66",x"cc"),
   895 => (x"d0",x"87",x"c7",x"03"),
   896 => (x"87",x"c2",x"02",x"66"),
   897 => (x"99",x"71",x"53",x"71"),
   898 => (x"c1",x"87",x"c2",x"02"),
   899 => (x"87",x"de",x"fd",x"84"),
   900 => (x"02",x"99",x"49",x"70"),
   901 => (x"ec",x"c0",x"87",x"cd"),
   902 => (x"87",x"c7",x"02",x"a9"),
   903 => (x"05",x"a9",x"fb",x"c0"),
   904 => (x"d0",x"87",x"d5",x"ff"),
   905 => (x"87",x"c3",x"02",x"66"),
   906 => (x"c0",x"7b",x"97",x"c0"),
   907 => (x"c4",x"05",x"a9",x"ec"),
   908 => (x"c5",x"4a",x"74",x"87"),
   909 => (x"c0",x"4a",x"74",x"87"),
   910 => (x"48",x"72",x"8a",x"0a"),
   911 => (x"4d",x"26",x"87",x"c2"),
   912 => (x"4b",x"26",x"4c",x"26"),
   913 => (x"fc",x"1e",x"4f",x"26"),
   914 => (x"49",x"70",x"87",x"e4"),
   915 => (x"aa",x"f0",x"c0",x"4a"),
   916 => (x"c0",x"87",x"c9",x"04"),
   917 => (x"c3",x"01",x"aa",x"f9"),
   918 => (x"8a",x"f0",x"c0",x"87"),
   919 => (x"04",x"aa",x"c1",x"c1"),
   920 => (x"da",x"c1",x"87",x"c9"),
   921 => (x"87",x"c3",x"01",x"aa"),
   922 => (x"72",x"8a",x"f7",x"c0"),
   923 => (x"0e",x"4f",x"26",x"48"),
   924 => (x"0e",x"5c",x"5b",x"5e"),
   925 => (x"d4",x"ff",x"4a",x"71"),
   926 => (x"c0",x"49",x"72",x"4c"),
   927 => (x"4b",x"70",x"87",x"e9"),
   928 => (x"87",x"c2",x"02",x"9b"),
   929 => (x"d0",x"ff",x"8b",x"c1"),
   930 => (x"c1",x"78",x"c5",x"48"),
   931 => (x"49",x"73",x"7c",x"d5"),
   932 => (x"e7",x"c1",x"31",x"c6"),
   933 => (x"4a",x"bf",x"97",x"c9"),
   934 => (x"70",x"b0",x"71",x"48"),
   935 => (x"48",x"d0",x"ff",x"7c"),
   936 => (x"48",x"73",x"78",x"c4"),
   937 => (x"0e",x"87",x"d9",x"fe"),
   938 => (x"5d",x"5c",x"5b",x"5e"),
   939 => (x"71",x"86",x"f4",x"0e"),
   940 => (x"48",x"a6",x"c4",x"4c"),
   941 => (x"a4",x"c8",x"78",x"c0"),
   942 => (x"bf",x"97",x"6e",x"7e"),
   943 => (x"a9",x"c1",x"c1",x"49"),
   944 => (x"c9",x"87",x"dd",x"05"),
   945 => (x"69",x"97",x"49",x"a4"),
   946 => (x"a9",x"d2",x"c1",x"49"),
   947 => (x"ca",x"87",x"d1",x"05"),
   948 => (x"69",x"97",x"49",x"a4"),
   949 => (x"a9",x"c3",x"c1",x"49"),
   950 => (x"df",x"87",x"c5",x"05"),
   951 => (x"87",x"e1",x"c2",x"48"),
   952 => (x"c0",x"87",x"eb",x"fa"),
   953 => (x"c6",x"fe",x"c0",x"4b"),
   954 => (x"c0",x"49",x"bf",x"97"),
   955 => (x"87",x"cf",x"04",x"a9"),
   956 => (x"c1",x"87",x"d0",x"fb"),
   957 => (x"c6",x"fe",x"c0",x"83"),
   958 => (x"ab",x"49",x"bf",x"97"),
   959 => (x"c0",x"87",x"f1",x"06"),
   960 => (x"bf",x"97",x"c6",x"fe"),
   961 => (x"f9",x"87",x"cf",x"02"),
   962 => (x"49",x"70",x"87",x"e4"),
   963 => (x"87",x"c6",x"02",x"99"),
   964 => (x"05",x"a9",x"ec",x"c0"),
   965 => (x"4b",x"c0",x"87",x"f1"),
   966 => (x"70",x"87",x"d3",x"f9"),
   967 => (x"87",x"ce",x"f9",x"4d"),
   968 => (x"f9",x"58",x"a6",x"cc"),
   969 => (x"4a",x"70",x"87",x"c8"),
   970 => (x"97",x"6e",x"83",x"c1"),
   971 => (x"02",x"ad",x"49",x"bf"),
   972 => (x"ff",x"c0",x"87",x"c7"),
   973 => (x"ea",x"c0",x"05",x"ad"),
   974 => (x"49",x"a4",x"c9",x"87"),
   975 => (x"c8",x"49",x"69",x"97"),
   976 => (x"c7",x"02",x"a9",x"66"),
   977 => (x"ff",x"c0",x"48",x"87"),
   978 => (x"87",x"d7",x"05",x"a8"),
   979 => (x"97",x"49",x"a4",x"ca"),
   980 => (x"02",x"aa",x"49",x"69"),
   981 => (x"ff",x"c0",x"87",x"c6"),
   982 => (x"87",x"c7",x"05",x"aa"),
   983 => (x"c1",x"48",x"a6",x"c4"),
   984 => (x"c0",x"87",x"d3",x"78"),
   985 => (x"c6",x"02",x"ad",x"ec"),
   986 => (x"ad",x"fb",x"c0",x"87"),
   987 => (x"c0",x"87",x"c7",x"05"),
   988 => (x"48",x"a6",x"c4",x"4b"),
   989 => (x"66",x"c4",x"78",x"c1"),
   990 => (x"87",x"dc",x"fe",x"02"),
   991 => (x"73",x"87",x"fb",x"f8"),
   992 => (x"fa",x"8e",x"f4",x"48"),
   993 => (x"0e",x"00",x"87",x"f8"),
   994 => (x"5d",x"5c",x"5b",x"5e"),
   995 => (x"71",x"86",x"f8",x"0e"),
   996 => (x"4b",x"d4",x"ff",x"4d"),
   997 => (x"f2",x"c2",x"1e",x"75"),
   998 => (x"df",x"ff",x"49",x"d8"),
   999 => (x"86",x"c4",x"87",x"e7"),
  1000 => (x"c4",x"02",x"98",x"70"),
  1001 => (x"e7",x"c1",x"87",x"fb"),
  1002 => (x"75",x"7e",x"bf",x"cb"),
  1003 => (x"87",x"ff",x"fa",x"49"),
  1004 => (x"c0",x"05",x"a8",x"de"),
  1005 => (x"49",x"75",x"87",x"eb"),
  1006 => (x"87",x"f9",x"f6",x"c0"),
  1007 => (x"db",x"02",x"98",x"70"),
  1008 => (x"fc",x"f6",x"c2",x"87"),
  1009 => (x"e1",x"c0",x"1e",x"bf"),
  1010 => (x"c8",x"f4",x"c0",x"49"),
  1011 => (x"c1",x"86",x"c4",x"87"),
  1012 => (x"c0",x"48",x"c9",x"e7"),
  1013 => (x"c8",x"f7",x"c2",x"50"),
  1014 => (x"87",x"eb",x"fe",x"49"),
  1015 => (x"c2",x"c4",x"48",x"c1"),
  1016 => (x"48",x"d0",x"ff",x"87"),
  1017 => (x"d6",x"c1",x"78",x"c5"),
  1018 => (x"75",x"4a",x"c0",x"7b"),
  1019 => (x"7b",x"11",x"49",x"a2"),
  1020 => (x"b7",x"cb",x"82",x"c1"),
  1021 => (x"87",x"f3",x"04",x"aa"),
  1022 => (x"ff",x"c3",x"4a",x"cc"),
  1023 => (x"c0",x"82",x"c1",x"7b"),
  1024 => (x"04",x"aa",x"b7",x"e0"),
  1025 => (x"d0",x"ff",x"87",x"f4"),
  1026 => (x"c3",x"78",x"c4",x"48"),
  1027 => (x"78",x"c5",x"7b",x"ff"),
  1028 => (x"c1",x"7b",x"d3",x"c1"),
  1029 => (x"6e",x"78",x"c4",x"7b"),
  1030 => (x"a8",x"b7",x"c0",x"48"),
  1031 => (x"87",x"f0",x"c2",x"06"),
  1032 => (x"bf",x"e0",x"f2",x"c2"),
  1033 => (x"74",x"48",x"6e",x"4c"),
  1034 => (x"74",x"7e",x"70",x"88"),
  1035 => (x"fd",x"c1",x"02",x"9c"),
  1036 => (x"e2",x"e5",x"c2",x"87"),
  1037 => (x"48",x"a6",x"c4",x"4d"),
  1038 => (x"8c",x"78",x"c0",x"c8"),
  1039 => (x"03",x"ac",x"b7",x"c0"),
  1040 => (x"c0",x"c8",x"87",x"c6"),
  1041 => (x"4c",x"c0",x"78",x"a4"),
  1042 => (x"97",x"d3",x"f2",x"c2"),
  1043 => (x"99",x"d0",x"49",x"bf"),
  1044 => (x"c0",x"87",x"d1",x"02"),
  1045 => (x"d8",x"f2",x"c2",x"1e"),
  1046 => (x"87",x"dc",x"e1",x"49"),
  1047 => (x"49",x"70",x"86",x"c4"),
  1048 => (x"87",x"ee",x"c0",x"4a"),
  1049 => (x"1e",x"e2",x"e5",x"c2"),
  1050 => (x"49",x"d8",x"f2",x"c2"),
  1051 => (x"c4",x"87",x"c9",x"e1"),
  1052 => (x"4a",x"49",x"70",x"86"),
  1053 => (x"c8",x"48",x"d0",x"ff"),
  1054 => (x"d4",x"c1",x"78",x"c5"),
  1055 => (x"c4",x"7b",x"15",x"7b"),
  1056 => (x"88",x"c1",x"48",x"66"),
  1057 => (x"70",x"58",x"a6",x"c8"),
  1058 => (x"f0",x"ff",x"05",x"98"),
  1059 => (x"48",x"d0",x"ff",x"87"),
  1060 => (x"9a",x"72",x"78",x"c4"),
  1061 => (x"c0",x"87",x"c5",x"05"),
  1062 => (x"87",x"c7",x"c1",x"48"),
  1063 => (x"f2",x"c2",x"1e",x"c1"),
  1064 => (x"de",x"ff",x"49",x"d8"),
  1065 => (x"86",x"c4",x"87",x"f8"),
  1066 => (x"fe",x"05",x"9c",x"74"),
  1067 => (x"48",x"6e",x"87",x"c3"),
  1068 => (x"06",x"a8",x"b7",x"c0"),
  1069 => (x"f2",x"c2",x"87",x"d1"),
  1070 => (x"78",x"c0",x"48",x"d8"),
  1071 => (x"78",x"c0",x"80",x"d0"),
  1072 => (x"f2",x"c2",x"80",x"f4"),
  1073 => (x"6e",x"78",x"bf",x"e4"),
  1074 => (x"a8",x"b7",x"c0",x"48"),
  1075 => (x"87",x"d0",x"fd",x"01"),
  1076 => (x"c5",x"48",x"d0",x"ff"),
  1077 => (x"7b",x"d3",x"c1",x"78"),
  1078 => (x"78",x"c4",x"7b",x"c0"),
  1079 => (x"c2",x"c0",x"48",x"c1"),
  1080 => (x"f8",x"48",x"c0",x"87"),
  1081 => (x"26",x"4d",x"26",x"8e"),
  1082 => (x"26",x"4b",x"26",x"4c"),
  1083 => (x"5b",x"5e",x"0e",x"4f"),
  1084 => (x"1e",x"0e",x"5d",x"5c"),
  1085 => (x"4c",x"c0",x"4b",x"71"),
  1086 => (x"c0",x"04",x"ab",x"4d"),
  1087 => (x"fa",x"c0",x"87",x"e8"),
  1088 => (x"9d",x"75",x"1e",x"e7"),
  1089 => (x"c0",x"87",x"c4",x"02"),
  1090 => (x"c1",x"87",x"c2",x"4a"),
  1091 => (x"e9",x"49",x"72",x"4a"),
  1092 => (x"86",x"c4",x"87",x"e2"),
  1093 => (x"84",x"c1",x"7e",x"70"),
  1094 => (x"87",x"c2",x"05",x"6e"),
  1095 => (x"85",x"c1",x"4c",x"73"),
  1096 => (x"ff",x"06",x"ac",x"73"),
  1097 => (x"48",x"6e",x"87",x"d8"),
  1098 => (x"87",x"f9",x"fe",x"26"),
  1099 => (x"c4",x"4a",x"71",x"1e"),
  1100 => (x"87",x"c5",x"05",x"66"),
  1101 => (x"ce",x"f9",x"49",x"72"),
  1102 => (x"0e",x"4f",x"26",x"87"),
  1103 => (x"5d",x"5c",x"5b",x"5e"),
  1104 => (x"4c",x"71",x"1e",x"0e"),
  1105 => (x"c2",x"91",x"de",x"49"),
  1106 => (x"71",x"4d",x"c0",x"f3"),
  1107 => (x"02",x"6d",x"97",x"85"),
  1108 => (x"c2",x"87",x"dc",x"c1"),
  1109 => (x"4a",x"bf",x"ec",x"f2"),
  1110 => (x"49",x"72",x"82",x"74"),
  1111 => (x"70",x"87",x"ce",x"fe"),
  1112 => (x"c0",x"02",x"6e",x"7e"),
  1113 => (x"f2",x"c2",x"87",x"f2"),
  1114 => (x"4a",x"6e",x"4b",x"f4"),
  1115 => (x"fc",x"fe",x"49",x"cb"),
  1116 => (x"4b",x"74",x"87",x"f6"),
  1117 => (x"e7",x"c1",x"93",x"cb"),
  1118 => (x"83",x"c4",x"83",x"dd"),
  1119 => (x"7b",x"f3",x"c6",x"c1"),
  1120 => (x"cb",x"c1",x"49",x"74"),
  1121 => (x"7b",x"75",x"87",x"d0"),
  1122 => (x"97",x"ca",x"e7",x"c1"),
  1123 => (x"c2",x"1e",x"49",x"bf"),
  1124 => (x"fe",x"49",x"f4",x"f2"),
  1125 => (x"86",x"c4",x"87",x"d6"),
  1126 => (x"ca",x"c1",x"49",x"74"),
  1127 => (x"49",x"c0",x"87",x"f8"),
  1128 => (x"87",x"d7",x"cc",x"c1"),
  1129 => (x"48",x"d4",x"f2",x"c2"),
  1130 => (x"49",x"c1",x"78",x"c0"),
  1131 => (x"26",x"87",x"d9",x"dd"),
  1132 => (x"4c",x"87",x"f2",x"fc"),
  1133 => (x"69",x"64",x"61",x"6f"),
  1134 => (x"2e",x"2e",x"67",x"6e"),
  1135 => (x"5e",x"0e",x"00",x"2e"),
  1136 => (x"71",x"0e",x"5c",x"5b"),
  1137 => (x"f2",x"c2",x"4a",x"4b"),
  1138 => (x"72",x"82",x"bf",x"ec"),
  1139 => (x"87",x"dd",x"fc",x"49"),
  1140 => (x"02",x"9c",x"4c",x"70"),
  1141 => (x"e5",x"49",x"87",x"c4"),
  1142 => (x"f2",x"c2",x"87",x"e2"),
  1143 => (x"78",x"c0",x"48",x"ec"),
  1144 => (x"e3",x"dc",x"49",x"c1"),
  1145 => (x"87",x"ff",x"fb",x"87"),
  1146 => (x"5c",x"5b",x"5e",x"0e"),
  1147 => (x"86",x"f4",x"0e",x"5d"),
  1148 => (x"4d",x"e2",x"e5",x"c2"),
  1149 => (x"a6",x"c4",x"4c",x"c0"),
  1150 => (x"c2",x"78",x"c0",x"48"),
  1151 => (x"49",x"bf",x"ec",x"f2"),
  1152 => (x"c1",x"06",x"a9",x"c0"),
  1153 => (x"e5",x"c2",x"87",x"c1"),
  1154 => (x"02",x"98",x"48",x"e2"),
  1155 => (x"c0",x"87",x"f8",x"c0"),
  1156 => (x"c8",x"1e",x"e7",x"fa"),
  1157 => (x"87",x"c7",x"02",x"66"),
  1158 => (x"c0",x"48",x"a6",x"c4"),
  1159 => (x"c4",x"87",x"c5",x"78"),
  1160 => (x"78",x"c1",x"48",x"a6"),
  1161 => (x"e5",x"49",x"66",x"c4"),
  1162 => (x"86",x"c4",x"87",x"ca"),
  1163 => (x"84",x"c1",x"4d",x"70"),
  1164 => (x"c1",x"48",x"66",x"c4"),
  1165 => (x"58",x"a6",x"c8",x"80"),
  1166 => (x"bf",x"ec",x"f2",x"c2"),
  1167 => (x"c6",x"03",x"ac",x"49"),
  1168 => (x"05",x"9d",x"75",x"87"),
  1169 => (x"c0",x"87",x"c8",x"ff"),
  1170 => (x"02",x"9d",x"75",x"4c"),
  1171 => (x"c0",x"87",x"e0",x"c3"),
  1172 => (x"c8",x"1e",x"e7",x"fa"),
  1173 => (x"87",x"c7",x"02",x"66"),
  1174 => (x"c0",x"48",x"a6",x"cc"),
  1175 => (x"cc",x"87",x"c5",x"78"),
  1176 => (x"78",x"c1",x"48",x"a6"),
  1177 => (x"e4",x"49",x"66",x"cc"),
  1178 => (x"86",x"c4",x"87",x"ca"),
  1179 => (x"02",x"6e",x"7e",x"70"),
  1180 => (x"6e",x"87",x"e9",x"c2"),
  1181 => (x"97",x"81",x"cb",x"49"),
  1182 => (x"99",x"d0",x"49",x"69"),
  1183 => (x"87",x"d6",x"c1",x"02"),
  1184 => (x"4a",x"fe",x"c6",x"c1"),
  1185 => (x"91",x"cb",x"49",x"74"),
  1186 => (x"81",x"dd",x"e7",x"c1"),
  1187 => (x"81",x"c8",x"79",x"72"),
  1188 => (x"74",x"51",x"ff",x"c3"),
  1189 => (x"c2",x"91",x"de",x"49"),
  1190 => (x"71",x"4d",x"c0",x"f3"),
  1191 => (x"97",x"c1",x"c2",x"85"),
  1192 => (x"49",x"a5",x"c1",x"7d"),
  1193 => (x"c2",x"51",x"e0",x"c0"),
  1194 => (x"bf",x"97",x"f2",x"ed"),
  1195 => (x"c1",x"87",x"d2",x"02"),
  1196 => (x"4b",x"a5",x"c2",x"84"),
  1197 => (x"4a",x"f2",x"ed",x"c2"),
  1198 => (x"f7",x"fe",x"49",x"db"),
  1199 => (x"db",x"c1",x"87",x"ea"),
  1200 => (x"49",x"a5",x"cd",x"87"),
  1201 => (x"84",x"c1",x"51",x"c0"),
  1202 => (x"6e",x"4b",x"a5",x"c2"),
  1203 => (x"fe",x"49",x"cb",x"4a"),
  1204 => (x"c1",x"87",x"d5",x"f7"),
  1205 => (x"c4",x"c1",x"87",x"c6"),
  1206 => (x"49",x"74",x"4a",x"fb"),
  1207 => (x"e7",x"c1",x"91",x"cb"),
  1208 => (x"79",x"72",x"81",x"dd"),
  1209 => (x"97",x"f2",x"ed",x"c2"),
  1210 => (x"87",x"d8",x"02",x"bf"),
  1211 => (x"91",x"de",x"49",x"74"),
  1212 => (x"f3",x"c2",x"84",x"c1"),
  1213 => (x"83",x"71",x"4b",x"c0"),
  1214 => (x"4a",x"f2",x"ed",x"c2"),
  1215 => (x"f6",x"fe",x"49",x"dd"),
  1216 => (x"87",x"d8",x"87",x"e6"),
  1217 => (x"93",x"de",x"4b",x"74"),
  1218 => (x"83",x"c0",x"f3",x"c2"),
  1219 => (x"c0",x"49",x"a3",x"cb"),
  1220 => (x"73",x"84",x"c1",x"51"),
  1221 => (x"49",x"cb",x"4a",x"6e"),
  1222 => (x"87",x"cc",x"f6",x"fe"),
  1223 => (x"c1",x"48",x"66",x"c4"),
  1224 => (x"58",x"a6",x"c8",x"80"),
  1225 => (x"c0",x"03",x"ac",x"c7"),
  1226 => (x"05",x"6e",x"87",x"c5"),
  1227 => (x"74",x"87",x"e0",x"fc"),
  1228 => (x"f6",x"8e",x"f4",x"48"),
  1229 => (x"73",x"1e",x"87",x"ef"),
  1230 => (x"49",x"4b",x"71",x"1e"),
  1231 => (x"e7",x"c1",x"91",x"cb"),
  1232 => (x"a1",x"c8",x"81",x"dd"),
  1233 => (x"c9",x"e7",x"c1",x"4a"),
  1234 => (x"c9",x"50",x"12",x"48"),
  1235 => (x"fe",x"c0",x"4a",x"a1"),
  1236 => (x"50",x"12",x"48",x"c6"),
  1237 => (x"e7",x"c1",x"81",x"ca"),
  1238 => (x"50",x"11",x"48",x"ca"),
  1239 => (x"97",x"ca",x"e7",x"c1"),
  1240 => (x"c0",x"1e",x"49",x"bf"),
  1241 => (x"87",x"c4",x"f7",x"49"),
  1242 => (x"48",x"d4",x"f2",x"c2"),
  1243 => (x"49",x"c1",x"78",x"de"),
  1244 => (x"26",x"87",x"d5",x"d6"),
  1245 => (x"1e",x"87",x"f2",x"f5"),
  1246 => (x"cb",x"49",x"4a",x"71"),
  1247 => (x"dd",x"e7",x"c1",x"91"),
  1248 => (x"11",x"81",x"c8",x"81"),
  1249 => (x"d8",x"f2",x"c2",x"48"),
  1250 => (x"ec",x"f2",x"c2",x"58"),
  1251 => (x"c1",x"78",x"c0",x"48"),
  1252 => (x"87",x"f4",x"d5",x"49"),
  1253 => (x"c0",x"1e",x"4f",x"26"),
  1254 => (x"de",x"c4",x"c1",x"49"),
  1255 => (x"1e",x"4f",x"26",x"87"),
  1256 => (x"d2",x"02",x"99",x"71"),
  1257 => (x"f2",x"e8",x"c1",x"87"),
  1258 => (x"f7",x"50",x"c0",x"48"),
  1259 => (x"f7",x"cd",x"c1",x"80"),
  1260 => (x"d6",x"e7",x"c1",x"40"),
  1261 => (x"c1",x"87",x"ce",x"78"),
  1262 => (x"c1",x"48",x"ee",x"e8"),
  1263 => (x"fc",x"78",x"cf",x"e7"),
  1264 => (x"d6",x"ce",x"c1",x"80"),
  1265 => (x"0e",x"4f",x"26",x"78"),
  1266 => (x"0e",x"5c",x"5b",x"5e"),
  1267 => (x"cb",x"4a",x"4c",x"71"),
  1268 => (x"dd",x"e7",x"c1",x"92"),
  1269 => (x"49",x"a2",x"c8",x"82"),
  1270 => (x"97",x"4b",x"a2",x"c9"),
  1271 => (x"97",x"1e",x"4b",x"6b"),
  1272 => (x"ca",x"1e",x"49",x"69"),
  1273 => (x"c0",x"49",x"12",x"82"),
  1274 => (x"c0",x"87",x"ca",x"e5"),
  1275 => (x"87",x"d8",x"d4",x"49"),
  1276 => (x"c1",x"c1",x"49",x"74"),
  1277 => (x"8e",x"f8",x"87",x"e0"),
  1278 => (x"1e",x"87",x"ec",x"f3"),
  1279 => (x"4b",x"71",x"1e",x"73"),
  1280 => (x"87",x"c3",x"ff",x"49"),
  1281 => (x"fe",x"fe",x"49",x"73"),
  1282 => (x"87",x"dd",x"f3",x"87"),
  1283 => (x"71",x"1e",x"73",x"1e"),
  1284 => (x"4a",x"a3",x"c6",x"4b"),
  1285 => (x"c1",x"87",x"db",x"02"),
  1286 => (x"87",x"d6",x"02",x"8a"),
  1287 => (x"da",x"c1",x"02",x"8a"),
  1288 => (x"c0",x"02",x"8a",x"87"),
  1289 => (x"02",x"8a",x"87",x"fc"),
  1290 => (x"8a",x"87",x"e1",x"c0"),
  1291 => (x"c1",x"87",x"cb",x"02"),
  1292 => (x"49",x"c7",x"87",x"db"),
  1293 => (x"c1",x"87",x"c0",x"fd"),
  1294 => (x"f2",x"c2",x"87",x"de"),
  1295 => (x"c1",x"02",x"bf",x"ec"),
  1296 => (x"c1",x"48",x"87",x"cb"),
  1297 => (x"f0",x"f2",x"c2",x"88"),
  1298 => (x"87",x"c1",x"c1",x"58"),
  1299 => (x"bf",x"f0",x"f2",x"c2"),
  1300 => (x"87",x"f9",x"c0",x"02"),
  1301 => (x"bf",x"ec",x"f2",x"c2"),
  1302 => (x"c2",x"80",x"c1",x"48"),
  1303 => (x"c0",x"58",x"f0",x"f2"),
  1304 => (x"f2",x"c2",x"87",x"eb"),
  1305 => (x"c6",x"49",x"bf",x"ec"),
  1306 => (x"f0",x"f2",x"c2",x"89"),
  1307 => (x"a9",x"b7",x"c0",x"59"),
  1308 => (x"c2",x"87",x"da",x"03"),
  1309 => (x"c0",x"48",x"ec",x"f2"),
  1310 => (x"c2",x"87",x"d2",x"78"),
  1311 => (x"02",x"bf",x"f0",x"f2"),
  1312 => (x"f2",x"c2",x"87",x"cb"),
  1313 => (x"c6",x"48",x"bf",x"ec"),
  1314 => (x"f0",x"f2",x"c2",x"80"),
  1315 => (x"d1",x"49",x"c0",x"58"),
  1316 => (x"49",x"73",x"87",x"f6"),
  1317 => (x"87",x"fe",x"fe",x"c0"),
  1318 => (x"1e",x"87",x"ce",x"f1"),
  1319 => (x"4b",x"71",x"1e",x"73"),
  1320 => (x"48",x"d4",x"f2",x"c2"),
  1321 => (x"49",x"c0",x"78",x"dd"),
  1322 => (x"73",x"87",x"dd",x"d1"),
  1323 => (x"e5",x"fe",x"c0",x"49"),
  1324 => (x"87",x"f5",x"f0",x"87"),
  1325 => (x"5c",x"5b",x"5e",x"0e"),
  1326 => (x"cc",x"ff",x"0e",x"5d"),
  1327 => (x"59",x"a6",x"d8",x"86"),
  1328 => (x"c0",x"48",x"a6",x"c8"),
  1329 => (x"c1",x"80",x"c4",x"78"),
  1330 => (x"c4",x"78",x"66",x"c8"),
  1331 => (x"c2",x"78",x"c1",x"80"),
  1332 => (x"c1",x"48",x"f0",x"f2"),
  1333 => (x"d4",x"f2",x"c2",x"78"),
  1334 => (x"a8",x"de",x"48",x"bf"),
  1335 => (x"f4",x"87",x"cb",x"05"),
  1336 => (x"49",x"70",x"87",x"c6"),
  1337 => (x"cf",x"59",x"a6",x"cc"),
  1338 => (x"e1",x"e2",x"87",x"d0"),
  1339 => (x"87",x"d3",x"e3",x"87"),
  1340 => (x"70",x"87",x"fb",x"e1"),
  1341 => (x"05",x"66",x"d4",x"4c"),
  1342 => (x"c1",x"87",x"fc",x"c1"),
  1343 => (x"c4",x"48",x"66",x"c4"),
  1344 => (x"c4",x"7e",x"70",x"80"),
  1345 => (x"bf",x"6e",x"48",x"a6"),
  1346 => (x"c1",x"1e",x"72",x"78"),
  1347 => (x"c8",x"48",x"ef",x"e3"),
  1348 => (x"a1",x"c8",x"49",x"66"),
  1349 => (x"71",x"41",x"20",x"4a"),
  1350 => (x"87",x"f9",x"05",x"aa"),
  1351 => (x"4a",x"26",x"51",x"10"),
  1352 => (x"48",x"66",x"c4",x"c1"),
  1353 => (x"78",x"f6",x"cc",x"c1"),
  1354 => (x"c7",x"49",x"bf",x"6e"),
  1355 => (x"c1",x"51",x"74",x"81"),
  1356 => (x"c8",x"49",x"66",x"c4"),
  1357 => (x"c1",x"51",x"c1",x"81"),
  1358 => (x"c9",x"49",x"66",x"c4"),
  1359 => (x"c1",x"51",x"c0",x"81"),
  1360 => (x"ca",x"49",x"66",x"c4"),
  1361 => (x"c0",x"51",x"c0",x"81"),
  1362 => (x"cf",x"02",x"ac",x"fb"),
  1363 => (x"d8",x"1e",x"c1",x"87"),
  1364 => (x"bf",x"66",x"c8",x"1e"),
  1365 => (x"e1",x"81",x"c8",x"49"),
  1366 => (x"86",x"c8",x"87",x"fd"),
  1367 => (x"48",x"66",x"c8",x"c1"),
  1368 => (x"c7",x"01",x"a8",x"c0"),
  1369 => (x"48",x"a6",x"c8",x"87"),
  1370 => (x"87",x"ce",x"78",x"c1"),
  1371 => (x"48",x"66",x"c8",x"c1"),
  1372 => (x"a6",x"d0",x"88",x"c1"),
  1373 => (x"e1",x"87",x"c3",x"58"),
  1374 => (x"a6",x"d8",x"87",x"c9"),
  1375 => (x"74",x"78",x"c2",x"48"),
  1376 => (x"f1",x"cc",x"02",x"9c"),
  1377 => (x"48",x"66",x"c8",x"87"),
  1378 => (x"a8",x"66",x"cc",x"c1"),
  1379 => (x"87",x"e6",x"cc",x"03"),
  1380 => (x"c0",x"48",x"a6",x"dc"),
  1381 => (x"c0",x"80",x"c4",x"78"),
  1382 => (x"d1",x"df",x"ff",x"78"),
  1383 => (x"d4",x"4c",x"70",x"87"),
  1384 => (x"a8",x"dd",x"48",x"66"),
  1385 => (x"c0",x"87",x"c7",x"05"),
  1386 => (x"d4",x"48",x"a6",x"e0"),
  1387 => (x"d0",x"c1",x"78",x"66"),
  1388 => (x"eb",x"c0",x"05",x"ac"),
  1389 => (x"f5",x"de",x"ff",x"87"),
  1390 => (x"f1",x"de",x"ff",x"87"),
  1391 => (x"c0",x"4c",x"70",x"87"),
  1392 => (x"c6",x"05",x"ac",x"ec"),
  1393 => (x"fa",x"df",x"ff",x"87"),
  1394 => (x"c1",x"4c",x"70",x"87"),
  1395 => (x"c8",x"05",x"ac",x"d0"),
  1396 => (x"48",x"66",x"d0",x"87"),
  1397 => (x"a6",x"d4",x"80",x"c1"),
  1398 => (x"ac",x"d0",x"c1",x"58"),
  1399 => (x"87",x"d5",x"ff",x"02"),
  1400 => (x"48",x"a6",x"e4",x"c0"),
  1401 => (x"c0",x"78",x"66",x"d4"),
  1402 => (x"c0",x"48",x"66",x"e0"),
  1403 => (x"05",x"a8",x"66",x"e4"),
  1404 => (x"c0",x"87",x"d5",x"ca"),
  1405 => (x"c0",x"48",x"a6",x"e8"),
  1406 => (x"80",x"dc",x"ff",x"78"),
  1407 => (x"4d",x"74",x"78",x"c0"),
  1408 => (x"02",x"8d",x"fb",x"c0"),
  1409 => (x"c9",x"87",x"db",x"c9"),
  1410 => (x"87",x"db",x"02",x"8d"),
  1411 => (x"c1",x"02",x"8d",x"c2"),
  1412 => (x"8d",x"c9",x"87",x"f7"),
  1413 => (x"87",x"d8",x"c4",x"02"),
  1414 => (x"c1",x"02",x"8d",x"c4"),
  1415 => (x"8d",x"c1",x"87",x"c1"),
  1416 => (x"87",x"cc",x"c4",x"02"),
  1417 => (x"c8",x"87",x"f5",x"c8"),
  1418 => (x"91",x"cb",x"49",x"66"),
  1419 => (x"81",x"66",x"c4",x"c1"),
  1420 => (x"6a",x"4a",x"a1",x"c4"),
  1421 => (x"c1",x"1e",x"71",x"7e"),
  1422 => (x"c4",x"48",x"fb",x"e3"),
  1423 => (x"a1",x"cc",x"49",x"66"),
  1424 => (x"71",x"41",x"20",x"4a"),
  1425 => (x"f8",x"ff",x"05",x"aa"),
  1426 => (x"26",x"51",x"10",x"87"),
  1427 => (x"db",x"d2",x"c1",x"49"),
  1428 => (x"d9",x"dc",x"ff",x"79"),
  1429 => (x"c4",x"4c",x"70",x"87"),
  1430 => (x"78",x"c1",x"48",x"a6"),
  1431 => (x"dc",x"87",x"c3",x"c8"),
  1432 => (x"f0",x"c0",x"48",x"a6"),
  1433 => (x"c5",x"dc",x"ff",x"78"),
  1434 => (x"c0",x"4c",x"70",x"87"),
  1435 => (x"c0",x"02",x"ac",x"ec"),
  1436 => (x"e0",x"c0",x"87",x"c4"),
  1437 => (x"ec",x"c0",x"5c",x"a6"),
  1438 => (x"87",x"cd",x"02",x"ac"),
  1439 => (x"87",x"ee",x"db",x"ff"),
  1440 => (x"ec",x"c0",x"4c",x"70"),
  1441 => (x"f3",x"ff",x"05",x"ac"),
  1442 => (x"ac",x"ec",x"c0",x"87"),
  1443 => (x"87",x"c4",x"c0",x"02"),
  1444 => (x"87",x"da",x"db",x"ff"),
  1445 => (x"1e",x"ca",x"1e",x"c0"),
  1446 => (x"cb",x"49",x"66",x"d0"),
  1447 => (x"66",x"cc",x"c1",x"91"),
  1448 => (x"cc",x"80",x"71",x"48"),
  1449 => (x"66",x"c8",x"58",x"a6"),
  1450 => (x"d0",x"80",x"c4",x"48"),
  1451 => (x"66",x"cc",x"58",x"a6"),
  1452 => (x"dc",x"ff",x"49",x"bf"),
  1453 => (x"1e",x"c1",x"87",x"e1"),
  1454 => (x"66",x"d4",x"1e",x"de"),
  1455 => (x"dc",x"ff",x"49",x"bf"),
  1456 => (x"86",x"d0",x"87",x"d5"),
  1457 => (x"09",x"c0",x"49",x"70"),
  1458 => (x"a6",x"f0",x"c0",x"89"),
  1459 => (x"66",x"ec",x"c0",x"59"),
  1460 => (x"06",x"a8",x"c0",x"48"),
  1461 => (x"c0",x"87",x"ee",x"c0"),
  1462 => (x"dd",x"48",x"66",x"ec"),
  1463 => (x"e4",x"c0",x"03",x"a8"),
  1464 => (x"bf",x"66",x"c4",x"87"),
  1465 => (x"66",x"ec",x"c0",x"49"),
  1466 => (x"51",x"e0",x"c0",x"81"),
  1467 => (x"49",x"66",x"ec",x"c0"),
  1468 => (x"66",x"c4",x"81",x"c1"),
  1469 => (x"c1",x"c2",x"81",x"bf"),
  1470 => (x"66",x"ec",x"c0",x"51"),
  1471 => (x"c4",x"81",x"c2",x"49"),
  1472 => (x"c0",x"81",x"bf",x"66"),
  1473 => (x"c1",x"48",x"6e",x"51"),
  1474 => (x"6e",x"78",x"f6",x"cc"),
  1475 => (x"d8",x"81",x"c8",x"49"),
  1476 => (x"49",x"6e",x"51",x"66"),
  1477 => (x"66",x"d0",x"81",x"c9"),
  1478 => (x"ca",x"49",x"6e",x"51"),
  1479 => (x"51",x"66",x"dc",x"81"),
  1480 => (x"c1",x"48",x"66",x"d8"),
  1481 => (x"58",x"a6",x"dc",x"80"),
  1482 => (x"c1",x"80",x"ec",x"48"),
  1483 => (x"87",x"f2",x"c4",x"78"),
  1484 => (x"87",x"d2",x"dc",x"ff"),
  1485 => (x"f0",x"c0",x"49",x"70"),
  1486 => (x"dc",x"ff",x"59",x"a6"),
  1487 => (x"49",x"70",x"87",x"c8"),
  1488 => (x"59",x"a6",x"e0",x"c0"),
  1489 => (x"c0",x"48",x"66",x"dc"),
  1490 => (x"c0",x"05",x"a8",x"ec"),
  1491 => (x"a6",x"dc",x"87",x"ca"),
  1492 => (x"66",x"ec",x"c0",x"48"),
  1493 => (x"87",x"c4",x"c0",x"78"),
  1494 => (x"87",x"d2",x"d8",x"ff"),
  1495 => (x"cb",x"49",x"66",x"c8"),
  1496 => (x"66",x"c4",x"c1",x"91"),
  1497 => (x"70",x"80",x"71",x"48"),
  1498 => (x"c8",x"4a",x"6e",x"7e"),
  1499 => (x"ca",x"49",x"6e",x"82"),
  1500 => (x"66",x"ec",x"c0",x"81"),
  1501 => (x"49",x"66",x"dc",x"51"),
  1502 => (x"ec",x"c0",x"81",x"c1"),
  1503 => (x"48",x"c1",x"89",x"66"),
  1504 => (x"49",x"70",x"30",x"71"),
  1505 => (x"97",x"71",x"89",x"c1"),
  1506 => (x"dc",x"f6",x"c2",x"7a"),
  1507 => (x"ec",x"c0",x"49",x"bf"),
  1508 => (x"6a",x"97",x"29",x"66"),
  1509 => (x"98",x"71",x"48",x"4a"),
  1510 => (x"58",x"a6",x"f4",x"c0"),
  1511 => (x"81",x"c4",x"49",x"6e"),
  1512 => (x"78",x"69",x"48",x"a6"),
  1513 => (x"48",x"66",x"e4",x"c0"),
  1514 => (x"a8",x"66",x"e0",x"c0"),
  1515 => (x"87",x"c8",x"c0",x"02"),
  1516 => (x"c0",x"48",x"a6",x"dc"),
  1517 => (x"87",x"c5",x"c0",x"78"),
  1518 => (x"c1",x"48",x"a6",x"dc"),
  1519 => (x"1e",x"66",x"dc",x"78"),
  1520 => (x"cc",x"1e",x"e0",x"c0"),
  1521 => (x"d8",x"ff",x"49",x"66"),
  1522 => (x"86",x"c8",x"87",x"cd"),
  1523 => (x"b7",x"c0",x"4c",x"70"),
  1524 => (x"db",x"c1",x"06",x"ac"),
  1525 => (x"48",x"66",x"c4",x"87"),
  1526 => (x"a6",x"c8",x"80",x"74"),
  1527 => (x"49",x"e0",x"c0",x"58"),
  1528 => (x"66",x"c4",x"89",x"74"),
  1529 => (x"f8",x"e3",x"c1",x"4b"),
  1530 => (x"e2",x"fe",x"71",x"4a"),
  1531 => (x"66",x"c4",x"87",x"fa"),
  1532 => (x"c8",x"80",x"c2",x"48"),
  1533 => (x"e8",x"c0",x"58",x"a6"),
  1534 => (x"80",x"c1",x"48",x"66"),
  1535 => (x"58",x"a6",x"ec",x"c0"),
  1536 => (x"49",x"66",x"f0",x"c0"),
  1537 => (x"a9",x"70",x"81",x"c1"),
  1538 => (x"87",x"c5",x"c0",x"02"),
  1539 => (x"c2",x"c0",x"4d",x"c0"),
  1540 => (x"75",x"4d",x"c1",x"87"),
  1541 => (x"49",x"a4",x"c2",x"1e"),
  1542 => (x"71",x"48",x"e0",x"c0"),
  1543 => (x"1e",x"49",x"70",x"88"),
  1544 => (x"ff",x"49",x"66",x"cc"),
  1545 => (x"c8",x"87",x"f0",x"d6"),
  1546 => (x"a8",x"b7",x"c0",x"86"),
  1547 => (x"87",x"c6",x"ff",x"01"),
  1548 => (x"02",x"66",x"e8",x"c0"),
  1549 => (x"6e",x"87",x"d1",x"c0"),
  1550 => (x"c0",x"81",x"c9",x"49"),
  1551 => (x"6e",x"51",x"66",x"e8"),
  1552 => (x"c7",x"cf",x"c1",x"48"),
  1553 => (x"87",x"cc",x"c0",x"78"),
  1554 => (x"81",x"c9",x"49",x"6e"),
  1555 => (x"48",x"6e",x"51",x"c2"),
  1556 => (x"78",x"fb",x"cf",x"c1"),
  1557 => (x"c1",x"48",x"a6",x"c4"),
  1558 => (x"87",x"c6",x"c0",x"78"),
  1559 => (x"87",x"e3",x"d5",x"ff"),
  1560 => (x"66",x"c4",x"4c",x"70"),
  1561 => (x"87",x"f5",x"c0",x"02"),
  1562 => (x"cc",x"48",x"66",x"c8"),
  1563 => (x"c0",x"04",x"a8",x"66"),
  1564 => (x"66",x"c8",x"87",x"cb"),
  1565 => (x"cc",x"80",x"c1",x"48"),
  1566 => (x"e0",x"c0",x"58",x"a6"),
  1567 => (x"48",x"66",x"cc",x"87"),
  1568 => (x"a6",x"d0",x"88",x"c1"),
  1569 => (x"87",x"d5",x"c0",x"58"),
  1570 => (x"05",x"ac",x"c6",x"c1"),
  1571 => (x"d8",x"87",x"c8",x"c0"),
  1572 => (x"80",x"c1",x"48",x"66"),
  1573 => (x"ff",x"58",x"a6",x"dc"),
  1574 => (x"70",x"87",x"e8",x"d4"),
  1575 => (x"48",x"66",x"d0",x"4c"),
  1576 => (x"a6",x"d4",x"80",x"c1"),
  1577 => (x"02",x"9c",x"74",x"58"),
  1578 => (x"c8",x"87",x"cb",x"c0"),
  1579 => (x"cc",x"c1",x"48",x"66"),
  1580 => (x"f3",x"04",x"a8",x"66"),
  1581 => (x"d4",x"ff",x"87",x"da"),
  1582 => (x"66",x"c8",x"87",x"c0"),
  1583 => (x"03",x"a8",x"c7",x"48"),
  1584 => (x"c2",x"87",x"e5",x"c0"),
  1585 => (x"c0",x"48",x"f0",x"f2"),
  1586 => (x"49",x"66",x"c8",x"78"),
  1587 => (x"c4",x"c1",x"91",x"cb"),
  1588 => (x"a1",x"c4",x"81",x"66"),
  1589 => (x"c0",x"4a",x"6a",x"4a"),
  1590 => (x"66",x"c8",x"79",x"52"),
  1591 => (x"cc",x"80",x"c1",x"48"),
  1592 => (x"a8",x"c7",x"58",x"a6"),
  1593 => (x"87",x"db",x"ff",x"04"),
  1594 => (x"ff",x"8e",x"cc",x"ff"),
  1595 => (x"4c",x"87",x"f6",x"df"),
  1596 => (x"20",x"64",x"61",x"6f"),
  1597 => (x"00",x"20",x"2e",x"2a"),
  1598 => (x"44",x"00",x"20",x"3a"),
  1599 => (x"53",x"20",x"50",x"49"),
  1600 => (x"63",x"74",x"69",x"77"),
  1601 => (x"00",x"73",x"65",x"68"),
  1602 => (x"71",x"1e",x"73",x"1e"),
  1603 => (x"c6",x"02",x"9b",x"4b"),
  1604 => (x"ec",x"f2",x"c2",x"87"),
  1605 => (x"c7",x"78",x"c0",x"48"),
  1606 => (x"ec",x"f2",x"c2",x"1e"),
  1607 => (x"c1",x"1e",x"49",x"bf"),
  1608 => (x"c2",x"1e",x"dd",x"e7"),
  1609 => (x"49",x"bf",x"d4",x"f2"),
  1610 => (x"cc",x"87",x"c9",x"ee"),
  1611 => (x"d4",x"f2",x"c2",x"86"),
  1612 => (x"ea",x"e9",x"49",x"bf"),
  1613 => (x"02",x"9b",x"73",x"87"),
  1614 => (x"e7",x"c1",x"87",x"c8"),
  1615 => (x"ed",x"c0",x"49",x"dd"),
  1616 => (x"de",x"ff",x"87",x"e6"),
  1617 => (x"c7",x"1e",x"87",x"e3"),
  1618 => (x"49",x"c1",x"87",x"cd"),
  1619 => (x"fe",x"87",x"f9",x"fe"),
  1620 => (x"70",x"87",x"e3",x"e5"),
  1621 => (x"87",x"cd",x"02",x"98"),
  1622 => (x"87",x"fc",x"ec",x"fe"),
  1623 => (x"c4",x"02",x"98",x"70"),
  1624 => (x"c2",x"4a",x"c1",x"87"),
  1625 => (x"72",x"4a",x"c0",x"87"),
  1626 => (x"87",x"ce",x"05",x"9a"),
  1627 => (x"e6",x"c1",x"1e",x"c0"),
  1628 => (x"f9",x"c0",x"49",x"db"),
  1629 => (x"86",x"c4",x"87",x"d0"),
  1630 => (x"fb",x"c0",x"87",x"fe"),
  1631 => (x"1e",x"c0",x"87",x"f3"),
  1632 => (x"49",x"e6",x"e6",x"c1"),
  1633 => (x"87",x"fe",x"f8",x"c0"),
  1634 => (x"fd",x"c0",x"1e",x"c0"),
  1635 => (x"49",x"70",x"87",x"f9"),
  1636 => (x"87",x"f2",x"f8",x"c0"),
  1637 => (x"f8",x"87",x"ff",x"c2"),
  1638 => (x"53",x"4f",x"26",x"8e"),
  1639 => (x"61",x"66",x"20",x"44"),
  1640 => (x"64",x"65",x"6c",x"69"),
  1641 => (x"6f",x"42",x"00",x"2e"),
  1642 => (x"6e",x"69",x"74",x"6f"),
  1643 => (x"2e",x"2e",x"2e",x"67"),
  1644 => (x"f2",x"c2",x"1e",x"00"),
  1645 => (x"78",x"c0",x"48",x"ec"),
  1646 => (x"48",x"d4",x"f2",x"c2"),
  1647 => (x"c5",x"fe",x"78",x"c0"),
  1648 => (x"e1",x"fd",x"c0",x"87"),
  1649 => (x"26",x"48",x"c0",x"87"),
  1650 => (x"01",x"00",x"00",x"4f"),
  1651 => (x"80",x"00",x"00",x"00"),
  1652 => (x"69",x"78",x"45",x"20"),
  1653 => (x"20",x"80",x"00",x"74"),
  1654 => (x"6b",x"63",x"61",x"42"),
  1655 => (x"00",x"13",x"77",x"00"),
  1656 => (x"00",x"2c",x"c0",x"00"),
  1657 => (x"00",x"00",x"00",x"00"),
  1658 => (x"00",x"00",x"13",x"77"),
  1659 => (x"00",x"00",x"2c",x"de"),
  1660 => (x"77",x"00",x"00",x"00"),
  1661 => (x"fc",x"00",x"00",x"13"),
  1662 => (x"00",x"00",x"00",x"2c"),
  1663 => (x"13",x"77",x"00",x"00"),
  1664 => (x"2d",x"1a",x"00",x"00"),
  1665 => (x"00",x"00",x"00",x"00"),
  1666 => (x"00",x"13",x"77",x"00"),
  1667 => (x"00",x"2d",x"38",x"00"),
  1668 => (x"00",x"00",x"00",x"00"),
  1669 => (x"00",x"00",x"13",x"77"),
  1670 => (x"00",x"00",x"2d",x"56"),
  1671 => (x"77",x"00",x"00",x"00"),
  1672 => (x"74",x"00",x"00",x"13"),
  1673 => (x"00",x"00",x"00",x"2d"),
  1674 => (x"13",x"77",x"00",x"00"),
  1675 => (x"00",x"00",x"00",x"00"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"00",x"14",x"0c",x"00"),
  1678 => (x"00",x"00",x"00",x"00"),
  1679 => (x"00",x"00",x"00",x"00"),
  1680 => (x"48",x"f0",x"fe",x"1e"),
  1681 => (x"09",x"cd",x"78",x"c0"),
  1682 => (x"4f",x"26",x"09",x"79"),
  1683 => (x"f0",x"fe",x"1e",x"1e"),
  1684 => (x"26",x"48",x"7e",x"bf"),
  1685 => (x"fe",x"1e",x"4f",x"26"),
  1686 => (x"78",x"c1",x"48",x"f0"),
  1687 => (x"fe",x"1e",x"4f",x"26"),
  1688 => (x"78",x"c0",x"48",x"f0"),
  1689 => (x"71",x"1e",x"4f",x"26"),
  1690 => (x"52",x"52",x"c0",x"4a"),
  1691 => (x"5e",x"0e",x"4f",x"26"),
  1692 => (x"0e",x"5d",x"5c",x"5b"),
  1693 => (x"4d",x"71",x"86",x"f4"),
  1694 => (x"c1",x"7e",x"6d",x"97"),
  1695 => (x"6c",x"97",x"4c",x"a5"),
  1696 => (x"58",x"a6",x"c8",x"48"),
  1697 => (x"66",x"c4",x"48",x"6e"),
  1698 => (x"87",x"c5",x"05",x"a8"),
  1699 => (x"e6",x"c0",x"48",x"ff"),
  1700 => (x"87",x"ca",x"ff",x"87"),
  1701 => (x"97",x"49",x"a5",x"c2"),
  1702 => (x"a3",x"71",x"4b",x"6c"),
  1703 => (x"4b",x"6b",x"97",x"4b"),
  1704 => (x"6e",x"7e",x"6c",x"97"),
  1705 => (x"c8",x"80",x"c1",x"48"),
  1706 => (x"98",x"c7",x"58",x"a6"),
  1707 => (x"70",x"58",x"a6",x"cc"),
  1708 => (x"e1",x"fe",x"7c",x"97"),
  1709 => (x"f4",x"48",x"73",x"87"),
  1710 => (x"26",x"4d",x"26",x"8e"),
  1711 => (x"26",x"4b",x"26",x"4c"),
  1712 => (x"5b",x"5e",x"0e",x"4f"),
  1713 => (x"86",x"f4",x"0e",x"5c"),
  1714 => (x"66",x"d8",x"4c",x"71"),
  1715 => (x"9a",x"ff",x"c3",x"4a"),
  1716 => (x"97",x"4b",x"a4",x"c2"),
  1717 => (x"a1",x"73",x"49",x"6c"),
  1718 => (x"97",x"51",x"72",x"49"),
  1719 => (x"48",x"6e",x"7e",x"6c"),
  1720 => (x"a6",x"c8",x"80",x"c1"),
  1721 => (x"cc",x"98",x"c7",x"58"),
  1722 => (x"54",x"70",x"58",x"a6"),
  1723 => (x"ca",x"ff",x"8e",x"f4"),
  1724 => (x"fd",x"1e",x"1e",x"87"),
  1725 => (x"bf",x"e0",x"87",x"e8"),
  1726 => (x"e0",x"c0",x"49",x"4a"),
  1727 => (x"cb",x"02",x"99",x"c0"),
  1728 => (x"c2",x"1e",x"72",x"87"),
  1729 => (x"fe",x"49",x"d2",x"f6"),
  1730 => (x"86",x"c4",x"87",x"f7"),
  1731 => (x"70",x"87",x"fd",x"fc"),
  1732 => (x"87",x"c2",x"fd",x"7e"),
  1733 => (x"1e",x"4f",x"26",x"26"),
  1734 => (x"49",x"d2",x"f6",x"c2"),
  1735 => (x"c1",x"87",x"c7",x"fd"),
  1736 => (x"fc",x"49",x"f1",x"eb"),
  1737 => (x"c7",x"c4",x"87",x"da"),
  1738 => (x"1e",x"4f",x"26",x"87"),
  1739 => (x"c8",x"48",x"d0",x"ff"),
  1740 => (x"d4",x"ff",x"78",x"e1"),
  1741 => (x"c4",x"78",x"c5",x"48"),
  1742 => (x"87",x"c3",x"02",x"66"),
  1743 => (x"c8",x"78",x"e0",x"c3"),
  1744 => (x"87",x"c6",x"02",x"66"),
  1745 => (x"c3",x"48",x"d4",x"ff"),
  1746 => (x"d4",x"ff",x"78",x"f0"),
  1747 => (x"ff",x"78",x"71",x"48"),
  1748 => (x"e1",x"c8",x"48",x"d0"),
  1749 => (x"78",x"e0",x"c0",x"78"),
  1750 => (x"5e",x"0e",x"4f",x"26"),
  1751 => (x"71",x"0e",x"5c",x"5b"),
  1752 => (x"d2",x"f6",x"c2",x"4c"),
  1753 => (x"87",x"c6",x"fc",x"49"),
  1754 => (x"b7",x"c0",x"4a",x"70"),
  1755 => (x"e2",x"c2",x"04",x"aa"),
  1756 => (x"aa",x"f0",x"c3",x"87"),
  1757 => (x"c1",x"87",x"c9",x"05"),
  1758 => (x"c1",x"48",x"df",x"f0"),
  1759 => (x"87",x"c3",x"c2",x"78"),
  1760 => (x"05",x"aa",x"e0",x"c3"),
  1761 => (x"f0",x"c1",x"87",x"c9"),
  1762 => (x"78",x"c1",x"48",x"e3"),
  1763 => (x"c1",x"87",x"f4",x"c1"),
  1764 => (x"02",x"bf",x"e3",x"f0"),
  1765 => (x"c0",x"c2",x"87",x"c6"),
  1766 => (x"87",x"c2",x"4b",x"a2"),
  1767 => (x"9c",x"74",x"4b",x"72"),
  1768 => (x"c1",x"87",x"d1",x"05"),
  1769 => (x"1e",x"bf",x"df",x"f0"),
  1770 => (x"bf",x"e3",x"f0",x"c1"),
  1771 => (x"fd",x"49",x"72",x"1e"),
  1772 => (x"86",x"c8",x"87",x"f9"),
  1773 => (x"bf",x"df",x"f0",x"c1"),
  1774 => (x"87",x"e0",x"c0",x"02"),
  1775 => (x"b7",x"c4",x"49",x"73"),
  1776 => (x"f1",x"c1",x"91",x"29"),
  1777 => (x"4a",x"73",x"81",x"ff"),
  1778 => (x"92",x"c2",x"9a",x"cf"),
  1779 => (x"30",x"72",x"48",x"c1"),
  1780 => (x"ba",x"ff",x"4a",x"70"),
  1781 => (x"98",x"69",x"48",x"72"),
  1782 => (x"87",x"db",x"79",x"70"),
  1783 => (x"b7",x"c4",x"49",x"73"),
  1784 => (x"f1",x"c1",x"91",x"29"),
  1785 => (x"4a",x"73",x"81",x"ff"),
  1786 => (x"92",x"c2",x"9a",x"cf"),
  1787 => (x"30",x"72",x"48",x"c3"),
  1788 => (x"69",x"48",x"4a",x"70"),
  1789 => (x"c1",x"79",x"70",x"b0"),
  1790 => (x"c0",x"48",x"e3",x"f0"),
  1791 => (x"df",x"f0",x"c1",x"78"),
  1792 => (x"c2",x"78",x"c0",x"48"),
  1793 => (x"f9",x"49",x"d2",x"f6"),
  1794 => (x"4a",x"70",x"87",x"e4"),
  1795 => (x"03",x"aa",x"b7",x"c0"),
  1796 => (x"c0",x"87",x"de",x"fd"),
  1797 => (x"26",x"87",x"c2",x"48"),
  1798 => (x"26",x"4c",x"26",x"4d"),
  1799 => (x"00",x"4f",x"26",x"4b"),
  1800 => (x"00",x"00",x"00",x"00"),
  1801 => (x"1e",x"00",x"00",x"00"),
  1802 => (x"fc",x"49",x"4a",x"71"),
  1803 => (x"4f",x"26",x"87",x"ec"),
  1804 => (x"72",x"4a",x"c0",x"1e"),
  1805 => (x"c1",x"91",x"c4",x"49"),
  1806 => (x"c0",x"81",x"ff",x"f1"),
  1807 => (x"d0",x"82",x"c1",x"79"),
  1808 => (x"ee",x"04",x"aa",x"b7"),
  1809 => (x"0e",x"4f",x"26",x"87"),
  1810 => (x"5d",x"5c",x"5b",x"5e"),
  1811 => (x"f8",x"4d",x"71",x"0e"),
  1812 => (x"4a",x"75",x"87",x"cc"),
  1813 => (x"92",x"2a",x"b7",x"c4"),
  1814 => (x"82",x"ff",x"f1",x"c1"),
  1815 => (x"9c",x"cf",x"4c",x"75"),
  1816 => (x"49",x"6a",x"94",x"c2"),
  1817 => (x"c3",x"2b",x"74",x"4b"),
  1818 => (x"74",x"48",x"c2",x"9b"),
  1819 => (x"ff",x"4c",x"70",x"30"),
  1820 => (x"71",x"48",x"74",x"bc"),
  1821 => (x"f7",x"7a",x"70",x"98"),
  1822 => (x"48",x"73",x"87",x"dc"),
  1823 => (x"00",x"87",x"d8",x"fe"),
  1824 => (x"00",x"00",x"00",x"00"),
  1825 => (x"00",x"00",x"00",x"00"),
  1826 => (x"00",x"00",x"00",x"00"),
  1827 => (x"00",x"00",x"00",x"00"),
  1828 => (x"00",x"00",x"00",x"00"),
  1829 => (x"00",x"00",x"00",x"00"),
  1830 => (x"00",x"00",x"00",x"00"),
  1831 => (x"00",x"00",x"00",x"00"),
  1832 => (x"00",x"00",x"00",x"00"),
  1833 => (x"00",x"00",x"00",x"00"),
  1834 => (x"00",x"00",x"00",x"00"),
  1835 => (x"00",x"00",x"00",x"00"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"00",x"00",x"00",x"00"),
  1838 => (x"00",x"00",x"00",x"00"),
  1839 => (x"1e",x"00",x"00",x"00"),
  1840 => (x"c8",x"48",x"d0",x"ff"),
  1841 => (x"48",x"71",x"78",x"e1"),
  1842 => (x"78",x"08",x"d4",x"ff"),
  1843 => (x"ff",x"48",x"66",x"c4"),
  1844 => (x"26",x"78",x"08",x"d4"),
  1845 => (x"4a",x"71",x"1e",x"4f"),
  1846 => (x"1e",x"49",x"66",x"c4"),
  1847 => (x"de",x"ff",x"49",x"72"),
  1848 => (x"48",x"d0",x"ff",x"87"),
  1849 => (x"26",x"78",x"e0",x"c0"),
  1850 => (x"73",x"1e",x"4f",x"26"),
  1851 => (x"c8",x"4b",x"71",x"1e"),
  1852 => (x"73",x"1e",x"49",x"66"),
  1853 => (x"a2",x"e0",x"c1",x"4a"),
  1854 => (x"87",x"d9",x"ff",x"49"),
  1855 => (x"26",x"87",x"c4",x"26"),
  1856 => (x"26",x"4c",x"26",x"4d"),
  1857 => (x"1e",x"4f",x"26",x"4b"),
  1858 => (x"c3",x"4a",x"d4",x"ff"),
  1859 => (x"d0",x"ff",x"7a",x"ff"),
  1860 => (x"78",x"e1",x"c0",x"48"),
  1861 => (x"f6",x"c2",x"7a",x"de"),
  1862 => (x"49",x"7a",x"bf",x"dc"),
  1863 => (x"70",x"28",x"c8",x"48"),
  1864 => (x"d0",x"48",x"71",x"7a"),
  1865 => (x"71",x"7a",x"70",x"28"),
  1866 => (x"70",x"28",x"d8",x"48"),
  1867 => (x"48",x"d0",x"ff",x"7a"),
  1868 => (x"26",x"78",x"e0",x"c0"),
  1869 => (x"5b",x"5e",x"0e",x"4f"),
  1870 => (x"71",x"0e",x"5d",x"5c"),
  1871 => (x"dc",x"f6",x"c2",x"4c"),
  1872 => (x"74",x"4b",x"4d",x"bf"),
  1873 => (x"9b",x"66",x"d0",x"2b"),
  1874 => (x"66",x"d4",x"83",x"c1"),
  1875 => (x"87",x"c2",x"04",x"ab"),
  1876 => (x"4a",x"74",x"4b",x"c0"),
  1877 => (x"72",x"49",x"66",x"d0"),
  1878 => (x"75",x"b9",x"ff",x"31"),
  1879 => (x"72",x"48",x"73",x"99"),
  1880 => (x"48",x"4a",x"70",x"30"),
  1881 => (x"f6",x"c2",x"b0",x"71"),
  1882 => (x"da",x"fe",x"58",x"e0"),
  1883 => (x"26",x"4d",x"26",x"87"),
  1884 => (x"26",x"4b",x"26",x"4c"),
  1885 => (x"5b",x"5e",x"0e",x"4f"),
  1886 => (x"1e",x"0e",x"5d",x"5c"),
  1887 => (x"f6",x"c2",x"4c",x"71"),
  1888 => (x"4a",x"c0",x"4b",x"e0"),
  1889 => (x"fe",x"49",x"f4",x"c0"),
  1890 => (x"74",x"87",x"ed",x"cc"),
  1891 => (x"e0",x"f6",x"c2",x"1e"),
  1892 => (x"f0",x"e7",x"fe",x"49"),
  1893 => (x"70",x"86",x"c4",x"87"),
  1894 => (x"c0",x"02",x"99",x"49"),
  1895 => (x"1e",x"c4",x"87",x"ea"),
  1896 => (x"c2",x"1e",x"4d",x"a6"),
  1897 => (x"fe",x"49",x"e0",x"f6"),
  1898 => (x"c8",x"87",x"c7",x"ef"),
  1899 => (x"02",x"98",x"70",x"86"),
  1900 => (x"4a",x"75",x"87",x"d6"),
  1901 => (x"49",x"fe",x"f7",x"c1"),
  1902 => (x"ca",x"fe",x"4b",x"c4"),
  1903 => (x"98",x"70",x"87",x"ec"),
  1904 => (x"c0",x"87",x"ca",x"02"),
  1905 => (x"87",x"ed",x"c0",x"48"),
  1906 => (x"e8",x"c0",x"48",x"c0"),
  1907 => (x"87",x"f3",x"c0",x"87"),
  1908 => (x"70",x"87",x"c4",x"c1"),
  1909 => (x"87",x"c8",x"02",x"98"),
  1910 => (x"70",x"87",x"fc",x"c0"),
  1911 => (x"87",x"f8",x"05",x"98"),
  1912 => (x"bf",x"c0",x"f7",x"c2"),
  1913 => (x"c2",x"87",x"cc",x"02"),
  1914 => (x"c2",x"48",x"dc",x"f6"),
  1915 => (x"78",x"bf",x"c0",x"f7"),
  1916 => (x"c1",x"87",x"d4",x"fc"),
  1917 => (x"4d",x"26",x"26",x"48"),
  1918 => (x"4b",x"26",x"4c",x"26"),
  1919 => (x"41",x"5b",x"4f",x"26"),
  1920 => (x"1e",x"00",x"43",x"52"),
  1921 => (x"f6",x"c2",x"1e",x"c0"),
  1922 => (x"eb",x"fe",x"49",x"e0"),
  1923 => (x"f6",x"c2",x"87",x"f9"),
  1924 => (x"78",x"c0",x"48",x"f8"),
  1925 => (x"0e",x"4f",x"26",x"26"),
  1926 => (x"5d",x"5c",x"5b",x"5e"),
  1927 => (x"c0",x"86",x"f4",x"0e"),
  1928 => (x"f8",x"f6",x"c2",x"7e"),
  1929 => (x"b7",x"c3",x"48",x"bf"),
  1930 => (x"87",x"d1",x"03",x"a8"),
  1931 => (x"bf",x"f8",x"f6",x"c2"),
  1932 => (x"c2",x"80",x"c1",x"48"),
  1933 => (x"c0",x"58",x"fc",x"f6"),
  1934 => (x"d9",x"c6",x"48",x"fb"),
  1935 => (x"e0",x"f6",x"c2",x"87"),
  1936 => (x"c1",x"f1",x"fe",x"49"),
  1937 => (x"c0",x"4c",x"70",x"87"),
  1938 => (x"c4",x"03",x"ac",x"b7"),
  1939 => (x"c5",x"c6",x"48",x"87"),
  1940 => (x"f8",x"f6",x"c2",x"87"),
  1941 => (x"8a",x"c3",x"4a",x"bf"),
  1942 => (x"c1",x"87",x"d8",x"02"),
  1943 => (x"c7",x"c5",x"02",x"8a"),
  1944 => (x"c2",x"02",x"8a",x"87"),
  1945 => (x"02",x"8a",x"87",x"f2"),
  1946 => (x"8a",x"87",x"cf",x"c1"),
  1947 => (x"87",x"de",x"c3",x"02"),
  1948 => (x"c0",x"87",x"d9",x"c5"),
  1949 => (x"5c",x"a6",x"c8",x"4d"),
  1950 => (x"92",x"c4",x"4a",x"75"),
  1951 => (x"82",x"f4",x"ff",x"c1"),
  1952 => (x"4c",x"f4",x"f6",x"c2"),
  1953 => (x"6c",x"97",x"84",x"75"),
  1954 => (x"c1",x"4b",x"49",x"4b"),
  1955 => (x"6a",x"7c",x"97",x"a3"),
  1956 => (x"cc",x"48",x"11",x"81"),
  1957 => (x"66",x"c4",x"58",x"a6"),
  1958 => (x"a8",x"66",x"c8",x"48"),
  1959 => (x"c0",x"87",x"c3",x"02"),
  1960 => (x"66",x"c8",x"7c",x"97"),
  1961 => (x"c2",x"87",x"c7",x"05"),
  1962 => (x"c4",x"48",x"f8",x"f6"),
  1963 => (x"85",x"c1",x"78",x"a5"),
  1964 => (x"04",x"ad",x"b7",x"c4"),
  1965 => (x"c4",x"87",x"c1",x"ff"),
  1966 => (x"f7",x"c2",x"87",x"d2"),
  1967 => (x"c8",x"48",x"bf",x"c4"),
  1968 => (x"cb",x"01",x"a8",x"b7"),
  1969 => (x"02",x"ac",x"ca",x"87"),
  1970 => (x"ac",x"cd",x"87",x"c6"),
  1971 => (x"87",x"f3",x"c0",x"05"),
  1972 => (x"bf",x"c4",x"f7",x"c2"),
  1973 => (x"ab",x"b7",x"c8",x"4b"),
  1974 => (x"c2",x"87",x"d2",x"03"),
  1975 => (x"73",x"49",x"c8",x"f7"),
  1976 => (x"51",x"e0",x"c0",x"81"),
  1977 => (x"b7",x"c8",x"83",x"c1"),
  1978 => (x"ee",x"ff",x"04",x"ab"),
  1979 => (x"d0",x"f7",x"c2",x"87"),
  1980 => (x"50",x"d2",x"c1",x"48"),
  1981 => (x"c1",x"50",x"cf",x"c1"),
  1982 => (x"50",x"c0",x"50",x"cd"),
  1983 => (x"78",x"c3",x"80",x"e4"),
  1984 => (x"c2",x"87",x"c9",x"c3"),
  1985 => (x"49",x"bf",x"c4",x"f7"),
  1986 => (x"c2",x"80",x"c1",x"48"),
  1987 => (x"48",x"58",x"c8",x"f7"),
  1988 => (x"74",x"81",x"a0",x"c4"),
  1989 => (x"87",x"f4",x"c2",x"51"),
  1990 => (x"ac",x"b7",x"f0",x"c0"),
  1991 => (x"c0",x"87",x"da",x"04"),
  1992 => (x"01",x"ac",x"b7",x"f9"),
  1993 => (x"f6",x"c2",x"87",x"d3"),
  1994 => (x"ca",x"49",x"bf",x"fc"),
  1995 => (x"c0",x"4a",x"74",x"91"),
  1996 => (x"f6",x"c2",x"8a",x"f0"),
  1997 => (x"a1",x"72",x"48",x"fc"),
  1998 => (x"02",x"ac",x"ca",x"78"),
  1999 => (x"cd",x"87",x"c6",x"c0"),
  2000 => (x"c7",x"c2",x"05",x"ac"),
  2001 => (x"f8",x"f6",x"c2",x"87"),
  2002 => (x"c1",x"78",x"c3",x"48"),
  2003 => (x"f0",x"c0",x"87",x"fe"),
  2004 => (x"db",x"04",x"ac",x"b7"),
  2005 => (x"b7",x"f9",x"c0",x"87"),
  2006 => (x"d3",x"c0",x"01",x"ac"),
  2007 => (x"c0",x"f7",x"c2",x"87"),
  2008 => (x"91",x"d0",x"49",x"bf"),
  2009 => (x"f0",x"c0",x"4a",x"74"),
  2010 => (x"c0",x"f7",x"c2",x"8a"),
  2011 => (x"78",x"a1",x"72",x"48"),
  2012 => (x"ac",x"b7",x"c1",x"c1"),
  2013 => (x"87",x"db",x"c0",x"04"),
  2014 => (x"ac",x"b7",x"c6",x"c1"),
  2015 => (x"87",x"d3",x"c0",x"01"),
  2016 => (x"bf",x"c0",x"f7",x"c2"),
  2017 => (x"74",x"91",x"d0",x"49"),
  2018 => (x"8a",x"f7",x"c0",x"4a"),
  2019 => (x"48",x"c0",x"f7",x"c2"),
  2020 => (x"ca",x"78",x"a1",x"72"),
  2021 => (x"c6",x"c0",x"02",x"ac"),
  2022 => (x"05",x"ac",x"cd",x"87"),
  2023 => (x"c2",x"87",x"ed",x"c0"),
  2024 => (x"c3",x"48",x"f8",x"f6"),
  2025 => (x"87",x"e4",x"c0",x"78"),
  2026 => (x"05",x"ac",x"e2",x"c0"),
  2027 => (x"c0",x"87",x"c6",x"c0"),
  2028 => (x"d7",x"c0",x"7e",x"fb"),
  2029 => (x"02",x"ac",x"ca",x"87"),
  2030 => (x"cd",x"87",x"c6",x"c0"),
  2031 => (x"c9",x"c0",x"05",x"ac"),
  2032 => (x"f8",x"f6",x"c2",x"87"),
  2033 => (x"c0",x"78",x"c3",x"48"),
  2034 => (x"7e",x"74",x"87",x"c2"),
  2035 => (x"d0",x"f9",x"02",x"6e"),
  2036 => (x"c3",x"48",x"6e",x"87"),
  2037 => (x"8e",x"f4",x"99",x"ff"),
  2038 => (x"43",x"87",x"db",x"f8"),
  2039 => (x"3d",x"46",x"4e",x"4f"),
  2040 => (x"44",x"4f",x"4d",x"00"),
  2041 => (x"4d",x"41",x"4e",x"00"),
  2042 => (x"45",x"44",x"00",x"45"),
  2043 => (x"4c",x"55",x"41",x"46"),
  2044 => (x"00",x"30",x"3d",x"54"),
  2045 => (x"00",x"00",x"1f",x"db"),
  2046 => (x"00",x"00",x"1f",x"e1"),
  2047 => (x"00",x"00",x"1f",x"e5"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

