library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"454d414e",
     1 => x"46454400",
     2 => x"544c5541",
     3 => x"f600303d",
     4 => x"fc00001f",
     5 => x"0000001f",
     6 => x"05000020",
     7 => x"1e000020",
     8 => x"c848d0ff",
     9 => x"487178c9",
    10 => x"7808d4ff",
    11 => x"711e4f26",
    12 => x"87eb494a",
    13 => x"c848d0ff",
    14 => x"1e4f2678",
    15 => x"4b711e73",
    16 => x"bff8f7c2",
    17 => x"c287c302",
    18 => x"d0ff87eb",
    19 => x"78c9c848",
    20 => x"e0c04973",
    21 => x"48d4ffb1",
    22 => x"f7c27871",
    23 => x"78c048ec",
    24 => x"c50266c8",
    25 => x"49ffc387",
    26 => x"49c087c2",
    27 => x"59f4f7c2",
    28 => x"c60266cc",
    29 => x"d5d5c587",
    30 => x"cf87c44a",
    31 => x"c24affff",
    32 => x"c25af8f7",
    33 => x"c148f8f7",
    34 => x"2687c478",
    35 => x"264c264d",
    36 => x"0e4f264b",
    37 => x"5d5c5b5e",
    38 => x"c24a710e",
    39 => x"4cbff4f7",
    40 => x"cb029a72",
    41 => x"91c84987",
    42 => x"4bf1c0c2",
    43 => x"87c48371",
    44 => x"4bf1c4c2",
    45 => x"49134dc0",
    46 => x"f7c29974",
    47 => x"ffb9bff0",
    48 => x"787148d4",
    49 => x"852cb7c1",
    50 => x"04adb7c8",
    51 => x"f7c287e8",
    52 => x"c848bfec",
    53 => x"f0f7c280",
    54 => x"87effe58",
    55 => x"711e731e",
    56 => x"9a4a134b",
    57 => x"7287cb02",
    58 => x"87e7fe49",
    59 => x"059a4a13",
    60 => x"dafe87f5",
    61 => x"f7c21e87",
    62 => x"c249bfec",
    63 => x"c148ecf7",
    64 => x"c0c478a1",
    65 => x"db03a9b7",
    66 => x"48d4ff87",
    67 => x"bff0f7c2",
    68 => x"ecf7c278",
    69 => x"f7c249bf",
    70 => x"a1c148ec",
    71 => x"b7c0c478",
    72 => x"87e504a9",
    73 => x"c848d0ff",
    74 => x"f8f7c278",
    75 => x"2678c048",
    76 => x"0000004f",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00005f5f",
    80 => x"03030000",
    81 => x"00030300",
    82 => x"7f7f1400",
    83 => x"147f7f14",
    84 => x"2e240000",
    85 => x"123a6b6b",
    86 => x"366a4c00",
    87 => x"32566c18",
    88 => x"4f7e3000",
    89 => x"683a7759",
    90 => x"04000040",
    91 => x"00000307",
    92 => x"1c000000",
    93 => x"0041633e",
    94 => x"41000000",
    95 => x"001c3e63",
    96 => x"3e2a0800",
    97 => x"2a3e1c1c",
    98 => x"08080008",
    99 => x"08083e3e",
   100 => x"80000000",
   101 => x"000060e0",
   102 => x"08080000",
   103 => x"08080808",
   104 => x"00000000",
   105 => x"00006060",
   106 => x"30604000",
   107 => x"03060c18",
   108 => x"7f3e0001",
   109 => x"3e7f4d59",
   110 => x"06040000",
   111 => x"00007f7f",
   112 => x"63420000",
   113 => x"464f5971",
   114 => x"63220000",
   115 => x"367f4949",
   116 => x"161c1800",
   117 => x"107f7f13",
   118 => x"67270000",
   119 => x"397d4545",
   120 => x"7e3c0000",
   121 => x"3079494b",
   122 => x"01010000",
   123 => x"070f7971",
   124 => x"7f360000",
   125 => x"367f4949",
   126 => x"4f060000",
   127 => x"1e3f6949",
   128 => x"00000000",
   129 => x"00006666",
   130 => x"80000000",
   131 => x"000066e6",
   132 => x"08080000",
   133 => x"22221414",
   134 => x"14140000",
   135 => x"14141414",
   136 => x"22220000",
   137 => x"08081414",
   138 => x"03020000",
   139 => x"060f5951",
   140 => x"417f3e00",
   141 => x"1e1f555d",
   142 => x"7f7e0000",
   143 => x"7e7f0909",
   144 => x"7f7f0000",
   145 => x"367f4949",
   146 => x"3e1c0000",
   147 => x"41414163",
   148 => x"7f7f0000",
   149 => x"1c3e6341",
   150 => x"7f7f0000",
   151 => x"41414949",
   152 => x"7f7f0000",
   153 => x"01010909",
   154 => x"7f3e0000",
   155 => x"7a7b4941",
   156 => x"7f7f0000",
   157 => x"7f7f0808",
   158 => x"41000000",
   159 => x"00417f7f",
   160 => x"60200000",
   161 => x"3f7f4040",
   162 => x"087f7f00",
   163 => x"4163361c",
   164 => x"7f7f0000",
   165 => x"40404040",
   166 => x"067f7f00",
   167 => x"7f7f060c",
   168 => x"067f7f00",
   169 => x"7f7f180c",
   170 => x"7f3e0000",
   171 => x"3e7f4141",
   172 => x"7f7f0000",
   173 => x"060f0909",
   174 => x"417f3e00",
   175 => x"407e7f61",
   176 => x"7f7f0000",
   177 => x"667f1909",
   178 => x"6f260000",
   179 => x"327b594d",
   180 => x"01010000",
   181 => x"01017f7f",
   182 => x"7f3f0000",
   183 => x"3f7f4040",
   184 => x"3f0f0000",
   185 => x"0f3f7070",
   186 => x"307f7f00",
   187 => x"7f7f3018",
   188 => x"36634100",
   189 => x"63361c1c",
   190 => x"06030141",
   191 => x"03067c7c",
   192 => x"59716101",
   193 => x"4143474d",
   194 => x"7f000000",
   195 => x"0041417f",
   196 => x"06030100",
   197 => x"6030180c",
   198 => x"41000040",
   199 => x"007f7f41",
   200 => x"060c0800",
   201 => x"080c0603",
   202 => x"80808000",
   203 => x"80808080",
   204 => x"00000000",
   205 => x"00040703",
   206 => x"74200000",
   207 => x"787c5454",
   208 => x"7f7f0000",
   209 => x"387c4444",
   210 => x"7c380000",
   211 => x"00444444",
   212 => x"7c380000",
   213 => x"7f7f4444",
   214 => x"7c380000",
   215 => x"185c5454",
   216 => x"7e040000",
   217 => x"0005057f",
   218 => x"bc180000",
   219 => x"7cfca4a4",
   220 => x"7f7f0000",
   221 => x"787c0404",
   222 => x"00000000",
   223 => x"00407d3d",
   224 => x"80800000",
   225 => x"007dfd80",
   226 => x"7f7f0000",
   227 => x"446c3810",
   228 => x"00000000",
   229 => x"00407f3f",
   230 => x"0c7c7c00",
   231 => x"787c0c18",
   232 => x"7c7c0000",
   233 => x"787c0404",
   234 => x"7c380000",
   235 => x"387c4444",
   236 => x"fcfc0000",
   237 => x"183c2424",
   238 => x"3c180000",
   239 => x"fcfc2424",
   240 => x"7c7c0000",
   241 => x"080c0404",
   242 => x"5c480000",
   243 => x"20745454",
   244 => x"3f040000",
   245 => x"0044447f",
   246 => x"7c3c0000",
   247 => x"7c7c4040",
   248 => x"3c1c0000",
   249 => x"1c3c6060",
   250 => x"607c3c00",
   251 => x"3c7c6030",
   252 => x"386c4400",
   253 => x"446c3810",
   254 => x"bc1c0000",
   255 => x"1c3c60e0",
   256 => x"64440000",
   257 => x"444c5c74",
   258 => x"08080000",
   259 => x"4141773e",
   260 => x"00000000",
   261 => x"00007f7f",
   262 => x"41410000",
   263 => x"08083e77",
   264 => x"01010200",
   265 => x"01020203",
   266 => x"7f7f7f00",
   267 => x"7f7f7f7f",
   268 => x"1c080800",
   269 => x"7f3e3e1c",
   270 => x"3e7f7f7f",
   271 => x"081c1c3e",
   272 => x"18100008",
   273 => x"10187c7c",
   274 => x"30100000",
   275 => x"10307c7c",
   276 => x"60301000",
   277 => x"061e7860",
   278 => x"3c664200",
   279 => x"42663c18",
   280 => x"6a387800",
   281 => x"386cc6c2",
   282 => x"00006000",
   283 => x"60000060",
   284 => x"5b5e0e00",
   285 => x"1e0e5d5c",
   286 => x"f8c24c71",
   287 => x"c04dbfc9",
   288 => x"741ec04b",
   289 => x"87c702ab",
   290 => x"c048a6c4",
   291 => x"c487c578",
   292 => x"78c148a6",
   293 => x"731e66c4",
   294 => x"87dfee49",
   295 => x"e0c086c8",
   296 => x"87efef49",
   297 => x"6a4aa5c4",
   298 => x"87f0f049",
   299 => x"cb87c6f1",
   300 => x"c883c185",
   301 => x"ff04abb7",
   302 => x"262687c7",
   303 => x"264c264d",
   304 => x"1e4f264b",
   305 => x"f8c24a71",
   306 => x"f8c25acd",
   307 => x"78c748cd",
   308 => x"87ddfe49",
   309 => x"731e4f26",
   310 => x"c04a711e",
   311 => x"d303aab7",
   312 => x"f6e0c287",
   313 => x"87c405bf",
   314 => x"87c24bc1",
   315 => x"e0c24bc0",
   316 => x"87c45bfa",
   317 => x"5afae0c2",
   318 => x"bff6e0c2",
   319 => x"c19ac14a",
   320 => x"ec49a2c0",
   321 => x"48fc87e8",
   322 => x"bff6e0c2",
   323 => x"87effe78",
   324 => x"c44a711e",
   325 => x"49721e66",
   326 => x"87dddfff",
   327 => x"1e4f2626",
   328 => x"bff6e0c2",
   329 => x"cddcff49",
   330 => x"c1f8c287",
   331 => x"78bfe848",
   332 => x"48fdf7c2",
   333 => x"c278bfec",
   334 => x"4abfc1f8",
   335 => x"99ffc349",
   336 => x"722ab7c8",
   337 => x"c2b07148",
   338 => x"2658c9f8",
   339 => x"5b5e0e4f",
   340 => x"710e5d5c",
   341 => x"87c7ff4b",
   342 => x"48fcf7c2",
   343 => x"497350c0",
   344 => x"87f2dbff",
   345 => x"c24c4970",
   346 => x"49eecb9c",
   347 => x"7087cfcb",
   348 => x"f7c24d49",
   349 => x"05bf97fc",
   350 => x"d087e4c1",
   351 => x"f8c24966",
   352 => x"0599bfc5",
   353 => x"66d487d7",
   354 => x"fdf7c249",
   355 => x"cc0599bf",
   356 => x"ff497387",
   357 => x"7087ffda",
   358 => x"c2c10298",
   359 => x"fd4cc187",
   360 => x"497587fd",
   361 => x"7087e3ca",
   362 => x"87c60298",
   363 => x"48fcf7c2",
   364 => x"f7c250c1",
   365 => x"05bf97fc",
   366 => x"c287e4c0",
   367 => x"49bfc5f8",
   368 => x"059966d0",
   369 => x"c287d6ff",
   370 => x"49bffdf7",
   371 => x"059966d4",
   372 => x"7387caff",
   373 => x"fdd9ff49",
   374 => x"05987087",
   375 => x"7487fefe",
   376 => x"87d7fb48",
   377 => x"5c5b5e0e",
   378 => x"86f40e5d",
   379 => x"ec4c4dc0",
   380 => x"a6c47ebf",
   381 => x"c9f8c248",
   382 => x"1ec178bf",
   383 => x"49c71ec0",
   384 => x"c887cafd",
   385 => x"02987086",
   386 => x"49ff87ce",
   387 => x"c187c7fb",
   388 => x"d9ff49da",
   389 => x"4dc187c0",
   390 => x"97fcf7c2",
   391 => x"87c302bf",
   392 => x"c287c0c9",
   393 => x"4bbfc1f8",
   394 => x"bff6e0c2",
   395 => x"87ebc005",
   396 => x"ff49fdc3",
   397 => x"c387dfd8",
   398 => x"d8ff49fa",
   399 => x"497387d8",
   400 => x"7199ffc3",
   401 => x"fb49c01e",
   402 => x"497387c6",
   403 => x"7129b7c8",
   404 => x"fa49c11e",
   405 => x"86c887fa",
   406 => x"c287c1c6",
   407 => x"4bbfc5f8",
   408 => x"87dd029b",
   409 => x"bff2e0c2",
   410 => x"87dec749",
   411 => x"c4059870",
   412 => x"d24bc087",
   413 => x"49e0c287",
   414 => x"c287c3c7",
   415 => x"c658f6e0",
   416 => x"f2e0c287",
   417 => x"7378c048",
   418 => x"0599c249",
   419 => x"ebc387ce",
   420 => x"c1d7ff49",
   421 => x"c2497087",
   422 => x"87c20299",
   423 => x"49734cfb",
   424 => x"ce0599c1",
   425 => x"49f4c387",
   426 => x"87ead6ff",
   427 => x"99c24970",
   428 => x"fa87c202",
   429 => x"c849734c",
   430 => x"87ce0599",
   431 => x"ff49f5c3",
   432 => x"7087d3d6",
   433 => x"0299c249",
   434 => x"f8c287d5",
   435 => x"ca02bfcd",
   436 => x"88c14887",
   437 => x"58d1f8c2",
   438 => x"ff87c2c0",
   439 => x"734dc14c",
   440 => x"0599c449",
   441 => x"f2c387ce",
   442 => x"e9d5ff49",
   443 => x"c2497087",
   444 => x"87dc0299",
   445 => x"bfcdf8c2",
   446 => x"b7c7487e",
   447 => x"cbc003a8",
   448 => x"c1486e87",
   449 => x"d1f8c280",
   450 => x"87c2c058",
   451 => x"4dc14cfe",
   452 => x"ff49fdc3",
   453 => x"7087ffd4",
   454 => x"0299c249",
   455 => x"c287d5c0",
   456 => x"02bfcdf8",
   457 => x"c287c9c0",
   458 => x"c048cdf8",
   459 => x"87c2c078",
   460 => x"4dc14cfd",
   461 => x"ff49fac3",
   462 => x"7087dbd4",
   463 => x"0299c249",
   464 => x"c287d9c0",
   465 => x"48bfcdf8",
   466 => x"03a8b7c7",
   467 => x"c287c9c0",
   468 => x"c748cdf8",
   469 => x"87c2c078",
   470 => x"4dc14cfc",
   471 => x"03acb7c0",
   472 => x"c487d1c0",
   473 => x"d8c14a66",
   474 => x"c0026a82",
   475 => x"4b6a87c6",
   476 => x"0f734974",
   477 => x"f0c31ec0",
   478 => x"49dac11e",
   479 => x"c887cef7",
   480 => x"02987086",
   481 => x"c887e2c0",
   482 => x"f8c248a6",
   483 => x"c878bfcd",
   484 => x"91cb4966",
   485 => x"714866c4",
   486 => x"6e7e7080",
   487 => x"c8c002bf",
   488 => x"4bbf6e87",
   489 => x"734966c8",
   490 => x"029d750f",
   491 => x"c287c8c0",
   492 => x"49bfcdf8",
   493 => x"c287faf2",
   494 => x"02bffae0",
   495 => x"4987ddc0",
   496 => x"7087c7c2",
   497 => x"d3c00298",
   498 => x"cdf8c287",
   499 => x"e0f249bf",
   500 => x"f449c087",
   501 => x"e0c287c0",
   502 => x"78c048fa",
   503 => x"daf38ef4",
   504 => x"5b5e0e87",
   505 => x"1e0e5d5c",
   506 => x"f8c24c71",
   507 => x"c149bfc9",
   508 => x"c14da1cd",
   509 => x"7e6981d1",
   510 => x"cf029c74",
   511 => x"4ba5c487",
   512 => x"f8c27b74",
   513 => x"f249bfc9",
   514 => x"7b6e87f9",
   515 => x"c4059c74",
   516 => x"c24bc087",
   517 => x"734bc187",
   518 => x"87faf249",
   519 => x"c70266d4",
   520 => x"87da4987",
   521 => x"87c24a70",
   522 => x"e0c24ac0",
   523 => x"f2265afe",
   524 => x"000087c9",
   525 => x"00000000",
   526 => x"00000000",
   527 => x"711e0000",
   528 => x"bfc8ff4a",
   529 => x"48a17249",
   530 => x"ff1e4f26",
   531 => x"fe89bfc8",
   532 => x"c0c0c0c0",
   533 => x"c401a9c0",
   534 => x"c24ac087",
   535 => x"724ac187",
   536 => x"1e4f2648",
   537 => x"bff1e2c2",
   538 => x"c2b9c149",
   539 => x"ff59f5e2",
   540 => x"ffc348d4",
   541 => x"48d0ff78",
   542 => x"ff78e1c0",
   543 => x"78c148d4",
   544 => x"787131c4",
   545 => x"c048d0ff",
   546 => x"4f2678e0",
   547 => x"e5e2c21e",
   548 => x"f0f2c21e",
   549 => x"f9fbfd49",
   550 => x"7086c487",
   551 => x"87c30298",
   552 => x"2687c0ff",
   553 => x"4b35314f",
   554 => x"20205a48",
   555 => x"47464320",
   556 => x"00000000",
   557 => x"5b5e0e00",
   558 => x"c20e5d5c",
   559 => x"4abffdf7",
   560 => x"bfdee4c2",
   561 => x"bc724c49",
   562 => x"c6ff4d71",
   563 => x"4bc087df",
   564 => x"99d04974",
   565 => x"87e7c002",
   566 => x"c848d0ff",
   567 => x"d4ff78e1",
   568 => x"7578c548",
   569 => x"0299d049",
   570 => x"f0c387c3",
   571 => x"cce5c278",
   572 => x"11817349",
   573 => x"08d4ff48",
   574 => x"48d0ff78",
   575 => x"c178e0c0",
   576 => x"c8832d2c",
   577 => x"c7ff04ab",
   578 => x"d8c5ff87",
   579 => x"dee4c287",
   580 => x"fdf7c248",
   581 => x"4d2678bf",
   582 => x"4b264c26",
   583 => x"00004f26",
   584 => x"c11e0000",
   585 => x"de48d0e7",
   586 => x"f5e4c250",
   587 => x"e2d9fe49",
   588 => x"2648c087",
   589 => x"4f544a4f",
   590 => x"55525455",
   591 => x"4352414e",
   592 => x"dff21e00",
   593 => x"87edfd87",
   594 => x"4f2687f8",
   595 => x"25261e16",
   596 => x"3e3d362e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
