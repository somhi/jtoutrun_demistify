
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"5c",x"a6",x"c8",x"87"),
     1 => (x"03",x"ac",x"b7",x"c0"),
     2 => (x"48",x"87",x"c4",x"c0"),
     3 => (x"c4",x"87",x"ca",x"c0"),
     4 => (x"c6",x"f9",x"02",x"66"),
     5 => (x"ff",x"c3",x"48",x"87"),
     6 => (x"f8",x"8e",x"f4",x"99"),
     7 => (x"4f",x"43",x"87",x"cf"),
     8 => (x"00",x"3d",x"46",x"4e"),
     9 => (x"00",x"44",x"4f",x"4d"),
    10 => (x"45",x"4d",x"41",x"4e"),
    11 => (x"46",x"45",x"44",x"00"),
    12 => (x"54",x"4c",x"55",x"41"),
    13 => (x"1e",x"00",x"30",x"3d"),
    14 => (x"24",x"00",x"00",x"20"),
    15 => (x"28",x"00",x"00",x"20"),
    16 => (x"2d",x"00",x"00",x"20"),
    17 => (x"1e",x"00",x"00",x"20"),
    18 => (x"c8",x"48",x"d0",x"ff"),
    19 => (x"48",x"71",x"78",x"c9"),
    20 => (x"78",x"08",x"d4",x"ff"),
    21 => (x"71",x"1e",x"4f",x"26"),
    22 => (x"87",x"eb",x"49",x"4a"),
    23 => (x"c8",x"48",x"d0",x"ff"),
    24 => (x"1e",x"4f",x"26",x"78"),
    25 => (x"4b",x"71",x"1e",x"73"),
    26 => (x"bf",x"e0",x"f8",x"c2"),
    27 => (x"c2",x"87",x"c3",x"02"),
    28 => (x"d0",x"ff",x"87",x"eb"),
    29 => (x"78",x"c9",x"c8",x"48"),
    30 => (x"e0",x"c0",x"49",x"73"),
    31 => (x"48",x"d4",x"ff",x"b1"),
    32 => (x"f8",x"c2",x"78",x"71"),
    33 => (x"78",x"c0",x"48",x"d4"),
    34 => (x"c5",x"02",x"66",x"c8"),
    35 => (x"49",x"ff",x"c3",x"87"),
    36 => (x"49",x"c0",x"87",x"c2"),
    37 => (x"59",x"dc",x"f8",x"c2"),
    38 => (x"c6",x"02",x"66",x"cc"),
    39 => (x"d5",x"d5",x"c5",x"87"),
    40 => (x"cf",x"87",x"c4",x"4a"),
    41 => (x"c2",x"4a",x"ff",x"ff"),
    42 => (x"c2",x"5a",x"e0",x"f8"),
    43 => (x"c1",x"48",x"e0",x"f8"),
    44 => (x"26",x"87",x"c4",x"78"),
    45 => (x"26",x"4c",x"26",x"4d"),
    46 => (x"0e",x"4f",x"26",x"4b"),
    47 => (x"5d",x"5c",x"5b",x"5e"),
    48 => (x"c2",x"4a",x"71",x"0e"),
    49 => (x"4c",x"bf",x"dc",x"f8"),
    50 => (x"cb",x"02",x"9a",x"72"),
    51 => (x"91",x"c8",x"49",x"87"),
    52 => (x"4b",x"d9",x"c1",x"c2"),
    53 => (x"87",x"c4",x"83",x"71"),
    54 => (x"4b",x"d9",x"c5",x"c2"),
    55 => (x"49",x"13",x"4d",x"c0"),
    56 => (x"f8",x"c2",x"99",x"74"),
    57 => (x"ff",x"b9",x"bf",x"d8"),
    58 => (x"78",x"71",x"48",x"d4"),
    59 => (x"85",x"2c",x"b7",x"c1"),
    60 => (x"04",x"ad",x"b7",x"c8"),
    61 => (x"f8",x"c2",x"87",x"e8"),
    62 => (x"c8",x"48",x"bf",x"d4"),
    63 => (x"d8",x"f8",x"c2",x"80"),
    64 => (x"87",x"ef",x"fe",x"58"),
    65 => (x"71",x"1e",x"73",x"1e"),
    66 => (x"9a",x"4a",x"13",x"4b"),
    67 => (x"72",x"87",x"cb",x"02"),
    68 => (x"87",x"e7",x"fe",x"49"),
    69 => (x"05",x"9a",x"4a",x"13"),
    70 => (x"da",x"fe",x"87",x"f5"),
    71 => (x"f8",x"c2",x"1e",x"87"),
    72 => (x"c2",x"49",x"bf",x"d4"),
    73 => (x"c1",x"48",x"d4",x"f8"),
    74 => (x"c0",x"c4",x"78",x"a1"),
    75 => (x"db",x"03",x"a9",x"b7"),
    76 => (x"48",x"d4",x"ff",x"87"),
    77 => (x"bf",x"d8",x"f8",x"c2"),
    78 => (x"d4",x"f8",x"c2",x"78"),
    79 => (x"f8",x"c2",x"49",x"bf"),
    80 => (x"a1",x"c1",x"48",x"d4"),
    81 => (x"b7",x"c0",x"c4",x"78"),
    82 => (x"87",x"e5",x"04",x"a9"),
    83 => (x"c8",x"48",x"d0",x"ff"),
    84 => (x"e0",x"f8",x"c2",x"78"),
    85 => (x"26",x"78",x"c0",x"48"),
    86 => (x"00",x"00",x"00",x"4f"),
    87 => (x"00",x"00",x"00",x"00"),
    88 => (x"00",x"00",x"00",x"00"),
    89 => (x"00",x"00",x"5f",x"5f"),
    90 => (x"03",x"03",x"00",x"00"),
    91 => (x"00",x"03",x"03",x"00"),
    92 => (x"7f",x"7f",x"14",x"00"),
    93 => (x"14",x"7f",x"7f",x"14"),
    94 => (x"2e",x"24",x"00",x"00"),
    95 => (x"12",x"3a",x"6b",x"6b"),
    96 => (x"36",x"6a",x"4c",x"00"),
    97 => (x"32",x"56",x"6c",x"18"),
    98 => (x"4f",x"7e",x"30",x"00"),
    99 => (x"68",x"3a",x"77",x"59"),
   100 => (x"04",x"00",x"00",x"40"),
   101 => (x"00",x"00",x"03",x"07"),
   102 => (x"1c",x"00",x"00",x"00"),
   103 => (x"00",x"41",x"63",x"3e"),
   104 => (x"41",x"00",x"00",x"00"),
   105 => (x"00",x"1c",x"3e",x"63"),
   106 => (x"3e",x"2a",x"08",x"00"),
   107 => (x"2a",x"3e",x"1c",x"1c"),
   108 => (x"08",x"08",x"00",x"08"),
   109 => (x"08",x"08",x"3e",x"3e"),
   110 => (x"80",x"00",x"00",x"00"),
   111 => (x"00",x"00",x"60",x"e0"),
   112 => (x"08",x"08",x"00",x"00"),
   113 => (x"08",x"08",x"08",x"08"),
   114 => (x"00",x"00",x"00",x"00"),
   115 => (x"00",x"00",x"60",x"60"),
   116 => (x"30",x"60",x"40",x"00"),
   117 => (x"03",x"06",x"0c",x"18"),
   118 => (x"7f",x"3e",x"00",x"01"),
   119 => (x"3e",x"7f",x"4d",x"59"),
   120 => (x"06",x"04",x"00",x"00"),
   121 => (x"00",x"00",x"7f",x"7f"),
   122 => (x"63",x"42",x"00",x"00"),
   123 => (x"46",x"4f",x"59",x"71"),
   124 => (x"63",x"22",x"00",x"00"),
   125 => (x"36",x"7f",x"49",x"49"),
   126 => (x"16",x"1c",x"18",x"00"),
   127 => (x"10",x"7f",x"7f",x"13"),
   128 => (x"67",x"27",x"00",x"00"),
   129 => (x"39",x"7d",x"45",x"45"),
   130 => (x"7e",x"3c",x"00",x"00"),
   131 => (x"30",x"79",x"49",x"4b"),
   132 => (x"01",x"01",x"00",x"00"),
   133 => (x"07",x"0f",x"79",x"71"),
   134 => (x"7f",x"36",x"00",x"00"),
   135 => (x"36",x"7f",x"49",x"49"),
   136 => (x"4f",x"06",x"00",x"00"),
   137 => (x"1e",x"3f",x"69",x"49"),
   138 => (x"00",x"00",x"00",x"00"),
   139 => (x"00",x"00",x"66",x"66"),
   140 => (x"80",x"00",x"00",x"00"),
   141 => (x"00",x"00",x"66",x"e6"),
   142 => (x"08",x"08",x"00",x"00"),
   143 => (x"22",x"22",x"14",x"14"),
   144 => (x"14",x"14",x"00",x"00"),
   145 => (x"14",x"14",x"14",x"14"),
   146 => (x"22",x"22",x"00",x"00"),
   147 => (x"08",x"08",x"14",x"14"),
   148 => (x"03",x"02",x"00",x"00"),
   149 => (x"06",x"0f",x"59",x"51"),
   150 => (x"41",x"7f",x"3e",x"00"),
   151 => (x"1e",x"1f",x"55",x"5d"),
   152 => (x"7f",x"7e",x"00",x"00"),
   153 => (x"7e",x"7f",x"09",x"09"),
   154 => (x"7f",x"7f",x"00",x"00"),
   155 => (x"36",x"7f",x"49",x"49"),
   156 => (x"3e",x"1c",x"00",x"00"),
   157 => (x"41",x"41",x"41",x"63"),
   158 => (x"7f",x"7f",x"00",x"00"),
   159 => (x"1c",x"3e",x"63",x"41"),
   160 => (x"7f",x"7f",x"00",x"00"),
   161 => (x"41",x"41",x"49",x"49"),
   162 => (x"7f",x"7f",x"00",x"00"),
   163 => (x"01",x"01",x"09",x"09"),
   164 => (x"7f",x"3e",x"00",x"00"),
   165 => (x"7a",x"7b",x"49",x"41"),
   166 => (x"7f",x"7f",x"00",x"00"),
   167 => (x"7f",x"7f",x"08",x"08"),
   168 => (x"41",x"00",x"00",x"00"),
   169 => (x"00",x"41",x"7f",x"7f"),
   170 => (x"60",x"20",x"00",x"00"),
   171 => (x"3f",x"7f",x"40",x"40"),
   172 => (x"08",x"7f",x"7f",x"00"),
   173 => (x"41",x"63",x"36",x"1c"),
   174 => (x"7f",x"7f",x"00",x"00"),
   175 => (x"40",x"40",x"40",x"40"),
   176 => (x"06",x"7f",x"7f",x"00"),
   177 => (x"7f",x"7f",x"06",x"0c"),
   178 => (x"06",x"7f",x"7f",x"00"),
   179 => (x"7f",x"7f",x"18",x"0c"),
   180 => (x"7f",x"3e",x"00",x"00"),
   181 => (x"3e",x"7f",x"41",x"41"),
   182 => (x"7f",x"7f",x"00",x"00"),
   183 => (x"06",x"0f",x"09",x"09"),
   184 => (x"41",x"7f",x"3e",x"00"),
   185 => (x"40",x"7e",x"7f",x"61"),
   186 => (x"7f",x"7f",x"00",x"00"),
   187 => (x"66",x"7f",x"19",x"09"),
   188 => (x"6f",x"26",x"00",x"00"),
   189 => (x"32",x"7b",x"59",x"4d"),
   190 => (x"01",x"01",x"00",x"00"),
   191 => (x"01",x"01",x"7f",x"7f"),
   192 => (x"7f",x"3f",x"00",x"00"),
   193 => (x"3f",x"7f",x"40",x"40"),
   194 => (x"3f",x"0f",x"00",x"00"),
   195 => (x"0f",x"3f",x"70",x"70"),
   196 => (x"30",x"7f",x"7f",x"00"),
   197 => (x"7f",x"7f",x"30",x"18"),
   198 => (x"36",x"63",x"41",x"00"),
   199 => (x"63",x"36",x"1c",x"1c"),
   200 => (x"06",x"03",x"01",x"41"),
   201 => (x"03",x"06",x"7c",x"7c"),
   202 => (x"59",x"71",x"61",x"01"),
   203 => (x"41",x"43",x"47",x"4d"),
   204 => (x"7f",x"00",x"00",x"00"),
   205 => (x"00",x"41",x"41",x"7f"),
   206 => (x"06",x"03",x"01",x"00"),
   207 => (x"60",x"30",x"18",x"0c"),
   208 => (x"41",x"00",x"00",x"40"),
   209 => (x"00",x"7f",x"7f",x"41"),
   210 => (x"06",x"0c",x"08",x"00"),
   211 => (x"08",x"0c",x"06",x"03"),
   212 => (x"80",x"80",x"80",x"00"),
   213 => (x"80",x"80",x"80",x"80"),
   214 => (x"00",x"00",x"00",x"00"),
   215 => (x"00",x"04",x"07",x"03"),
   216 => (x"74",x"20",x"00",x"00"),
   217 => (x"78",x"7c",x"54",x"54"),
   218 => (x"7f",x"7f",x"00",x"00"),
   219 => (x"38",x"7c",x"44",x"44"),
   220 => (x"7c",x"38",x"00",x"00"),
   221 => (x"00",x"44",x"44",x"44"),
   222 => (x"7c",x"38",x"00",x"00"),
   223 => (x"7f",x"7f",x"44",x"44"),
   224 => (x"7c",x"38",x"00",x"00"),
   225 => (x"18",x"5c",x"54",x"54"),
   226 => (x"7e",x"04",x"00",x"00"),
   227 => (x"00",x"05",x"05",x"7f"),
   228 => (x"bc",x"18",x"00",x"00"),
   229 => (x"7c",x"fc",x"a4",x"a4"),
   230 => (x"7f",x"7f",x"00",x"00"),
   231 => (x"78",x"7c",x"04",x"04"),
   232 => (x"00",x"00",x"00",x"00"),
   233 => (x"00",x"40",x"7d",x"3d"),
   234 => (x"80",x"80",x"00",x"00"),
   235 => (x"00",x"7d",x"fd",x"80"),
   236 => (x"7f",x"7f",x"00",x"00"),
   237 => (x"44",x"6c",x"38",x"10"),
   238 => (x"00",x"00",x"00",x"00"),
   239 => (x"00",x"40",x"7f",x"3f"),
   240 => (x"0c",x"7c",x"7c",x"00"),
   241 => (x"78",x"7c",x"0c",x"18"),
   242 => (x"7c",x"7c",x"00",x"00"),
   243 => (x"78",x"7c",x"04",x"04"),
   244 => (x"7c",x"38",x"00",x"00"),
   245 => (x"38",x"7c",x"44",x"44"),
   246 => (x"fc",x"fc",x"00",x"00"),
   247 => (x"18",x"3c",x"24",x"24"),
   248 => (x"3c",x"18",x"00",x"00"),
   249 => (x"fc",x"fc",x"24",x"24"),
   250 => (x"7c",x"7c",x"00",x"00"),
   251 => (x"08",x"0c",x"04",x"04"),
   252 => (x"5c",x"48",x"00",x"00"),
   253 => (x"20",x"74",x"54",x"54"),
   254 => (x"3f",x"04",x"00",x"00"),
   255 => (x"00",x"44",x"44",x"7f"),
   256 => (x"7c",x"3c",x"00",x"00"),
   257 => (x"7c",x"7c",x"40",x"40"),
   258 => (x"3c",x"1c",x"00",x"00"),
   259 => (x"1c",x"3c",x"60",x"60"),
   260 => (x"60",x"7c",x"3c",x"00"),
   261 => (x"3c",x"7c",x"60",x"30"),
   262 => (x"38",x"6c",x"44",x"00"),
   263 => (x"44",x"6c",x"38",x"10"),
   264 => (x"bc",x"1c",x"00",x"00"),
   265 => (x"1c",x"3c",x"60",x"e0"),
   266 => (x"64",x"44",x"00",x"00"),
   267 => (x"44",x"4c",x"5c",x"74"),
   268 => (x"08",x"08",x"00",x"00"),
   269 => (x"41",x"41",x"77",x"3e"),
   270 => (x"00",x"00",x"00",x"00"),
   271 => (x"00",x"00",x"7f",x"7f"),
   272 => (x"41",x"41",x"00",x"00"),
   273 => (x"08",x"08",x"3e",x"77"),
   274 => (x"01",x"01",x"02",x"00"),
   275 => (x"01",x"02",x"02",x"03"),
   276 => (x"7f",x"7f",x"7f",x"00"),
   277 => (x"7f",x"7f",x"7f",x"7f"),
   278 => (x"1c",x"08",x"08",x"00"),
   279 => (x"7f",x"3e",x"3e",x"1c"),
   280 => (x"3e",x"7f",x"7f",x"7f"),
   281 => (x"08",x"1c",x"1c",x"3e"),
   282 => (x"18",x"10",x"00",x"08"),
   283 => (x"10",x"18",x"7c",x"7c"),
   284 => (x"30",x"10",x"00",x"00"),
   285 => (x"10",x"30",x"7c",x"7c"),
   286 => (x"60",x"30",x"10",x"00"),
   287 => (x"06",x"1e",x"78",x"60"),
   288 => (x"3c",x"66",x"42",x"00"),
   289 => (x"42",x"66",x"3c",x"18"),
   290 => (x"6a",x"38",x"78",x"00"),
   291 => (x"38",x"6c",x"c6",x"c2"),
   292 => (x"00",x"00",x"60",x"00"),
   293 => (x"60",x"00",x"00",x"60"),
   294 => (x"5b",x"5e",x"0e",x"00"),
   295 => (x"1e",x"0e",x"5d",x"5c"),
   296 => (x"f8",x"c2",x"4c",x"71"),
   297 => (x"c0",x"4d",x"bf",x"f1"),
   298 => (x"74",x"1e",x"c0",x"4b"),
   299 => (x"87",x"c7",x"02",x"ab"),
   300 => (x"c0",x"48",x"a6",x"c4"),
   301 => (x"c4",x"87",x"c5",x"78"),
   302 => (x"78",x"c1",x"48",x"a6"),
   303 => (x"73",x"1e",x"66",x"c4"),
   304 => (x"87",x"df",x"ee",x"49"),
   305 => (x"e0",x"c0",x"86",x"c8"),
   306 => (x"87",x"ef",x"ef",x"49"),
   307 => (x"6a",x"4a",x"a5",x"c4"),
   308 => (x"87",x"f0",x"f0",x"49"),
   309 => (x"cb",x"87",x"c6",x"f1"),
   310 => (x"c8",x"83",x"c1",x"85"),
   311 => (x"ff",x"04",x"ab",x"b7"),
   312 => (x"26",x"26",x"87",x"c7"),
   313 => (x"26",x"4c",x"26",x"4d"),
   314 => (x"1e",x"4f",x"26",x"4b"),
   315 => (x"f8",x"c2",x"4a",x"71"),
   316 => (x"f8",x"c2",x"5a",x"f5"),
   317 => (x"78",x"c7",x"48",x"f5"),
   318 => (x"87",x"dd",x"fe",x"49"),
   319 => (x"73",x"1e",x"4f",x"26"),
   320 => (x"c0",x"4a",x"71",x"1e"),
   321 => (x"d3",x"03",x"aa",x"b7"),
   322 => (x"de",x"e1",x"c2",x"87"),
   323 => (x"87",x"c4",x"05",x"bf"),
   324 => (x"87",x"c2",x"4b",x"c1"),
   325 => (x"e1",x"c2",x"4b",x"c0"),
   326 => (x"87",x"c4",x"5b",x"e2"),
   327 => (x"5a",x"e2",x"e1",x"c2"),
   328 => (x"bf",x"de",x"e1",x"c2"),
   329 => (x"c1",x"9a",x"c1",x"4a"),
   330 => (x"ec",x"49",x"a2",x"c0"),
   331 => (x"48",x"fc",x"87",x"e8"),
   332 => (x"bf",x"de",x"e1",x"c2"),
   333 => (x"87",x"ef",x"fe",x"78"),
   334 => (x"c4",x"4a",x"71",x"1e"),
   335 => (x"49",x"72",x"1e",x"66"),
   336 => (x"87",x"d2",x"df",x"ff"),
   337 => (x"1e",x"4f",x"26",x"26"),
   338 => (x"bf",x"de",x"e1",x"c2"),
   339 => (x"e5",x"db",x"ff",x"49"),
   340 => (x"e9",x"f8",x"c2",x"87"),
   341 => (x"78",x"bf",x"e8",x"48"),
   342 => (x"48",x"e5",x"f8",x"c2"),
   343 => (x"c2",x"78",x"bf",x"ec"),
   344 => (x"4a",x"bf",x"e9",x"f8"),
   345 => (x"99",x"ff",x"c3",x"49"),
   346 => (x"72",x"2a",x"b7",x"c8"),
   347 => (x"c2",x"b0",x"71",x"48"),
   348 => (x"26",x"58",x"f1",x"f8"),
   349 => (x"5b",x"5e",x"0e",x"4f"),
   350 => (x"71",x"0e",x"5d",x"5c"),
   351 => (x"87",x"c7",x"ff",x"4b"),
   352 => (x"48",x"e4",x"f8",x"c2"),
   353 => (x"49",x"73",x"50",x"c0"),
   354 => (x"87",x"ca",x"db",x"ff"),
   355 => (x"c2",x"4c",x"49",x"70"),
   356 => (x"49",x"ee",x"cb",x"9c"),
   357 => (x"70",x"87",x"cf",x"cb"),
   358 => (x"f8",x"c2",x"4d",x"49"),
   359 => (x"05",x"bf",x"97",x"e4"),
   360 => (x"d0",x"87",x"e4",x"c1"),
   361 => (x"f8",x"c2",x"49",x"66"),
   362 => (x"05",x"99",x"bf",x"ed"),
   363 => (x"66",x"d4",x"87",x"d7"),
   364 => (x"e5",x"f8",x"c2",x"49"),
   365 => (x"cc",x"05",x"99",x"bf"),
   366 => (x"ff",x"49",x"73",x"87"),
   367 => (x"70",x"87",x"d7",x"da"),
   368 => (x"c2",x"c1",x"02",x"98"),
   369 => (x"fd",x"4c",x"c1",x"87"),
   370 => (x"49",x"75",x"87",x"fd"),
   371 => (x"70",x"87",x"e3",x"ca"),
   372 => (x"87",x"c6",x"02",x"98"),
   373 => (x"48",x"e4",x"f8",x"c2"),
   374 => (x"f8",x"c2",x"50",x"c1"),
   375 => (x"05",x"bf",x"97",x"e4"),
   376 => (x"c2",x"87",x"e4",x"c0"),
   377 => (x"49",x"bf",x"ed",x"f8"),
   378 => (x"05",x"99",x"66",x"d0"),
   379 => (x"c2",x"87",x"d6",x"ff"),
   380 => (x"49",x"bf",x"e5",x"f8"),
   381 => (x"05",x"99",x"66",x"d4"),
   382 => (x"73",x"87",x"ca",x"ff"),
   383 => (x"d5",x"d9",x"ff",x"49"),
   384 => (x"05",x"98",x"70",x"87"),
   385 => (x"74",x"87",x"fe",x"fe"),
   386 => (x"87",x"d7",x"fb",x"48"),
   387 => (x"5c",x"5b",x"5e",x"0e"),
   388 => (x"86",x"f4",x"0e",x"5d"),
   389 => (x"ec",x"4c",x"4d",x"c0"),
   390 => (x"a6",x"c4",x"7e",x"bf"),
   391 => (x"f1",x"f8",x"c2",x"48"),
   392 => (x"1e",x"c1",x"78",x"bf"),
   393 => (x"49",x"c7",x"1e",x"c0"),
   394 => (x"c8",x"87",x"ca",x"fd"),
   395 => (x"02",x"98",x"70",x"86"),
   396 => (x"49",x"ff",x"87",x"ce"),
   397 => (x"c1",x"87",x"c7",x"fb"),
   398 => (x"d8",x"ff",x"49",x"da"),
   399 => (x"4d",x"c1",x"87",x"d8"),
   400 => (x"97",x"e4",x"f8",x"c2"),
   401 => (x"87",x"c3",x"02",x"bf"),
   402 => (x"c2",x"87",x"c0",x"c9"),
   403 => (x"4b",x"bf",x"e9",x"f8"),
   404 => (x"bf",x"de",x"e1",x"c2"),
   405 => (x"87",x"eb",x"c0",x"05"),
   406 => (x"ff",x"49",x"fd",x"c3"),
   407 => (x"c3",x"87",x"f7",x"d7"),
   408 => (x"d7",x"ff",x"49",x"fa"),
   409 => (x"49",x"73",x"87",x"f0"),
   410 => (x"71",x"99",x"ff",x"c3"),
   411 => (x"fb",x"49",x"c0",x"1e"),
   412 => (x"49",x"73",x"87",x"c6"),
   413 => (x"71",x"29",x"b7",x"c8"),
   414 => (x"fa",x"49",x"c1",x"1e"),
   415 => (x"86",x"c8",x"87",x"fa"),
   416 => (x"c2",x"87",x"c1",x"c6"),
   417 => (x"4b",x"bf",x"ed",x"f8"),
   418 => (x"87",x"dd",x"02",x"9b"),
   419 => (x"bf",x"da",x"e1",x"c2"),
   420 => (x"87",x"de",x"c7",x"49"),
   421 => (x"c4",x"05",x"98",x"70"),
   422 => (x"d2",x"4b",x"c0",x"87"),
   423 => (x"49",x"e0",x"c2",x"87"),
   424 => (x"c2",x"87",x"c3",x"c7"),
   425 => (x"c6",x"58",x"de",x"e1"),
   426 => (x"da",x"e1",x"c2",x"87"),
   427 => (x"73",x"78",x"c0",x"48"),
   428 => (x"05",x"99",x"c2",x"49"),
   429 => (x"eb",x"c3",x"87",x"ce"),
   430 => (x"d9",x"d6",x"ff",x"49"),
   431 => (x"c2",x"49",x"70",x"87"),
   432 => (x"87",x"c2",x"02",x"99"),
   433 => (x"49",x"73",x"4c",x"fb"),
   434 => (x"ce",x"05",x"99",x"c1"),
   435 => (x"49",x"f4",x"c3",x"87"),
   436 => (x"87",x"c2",x"d6",x"ff"),
   437 => (x"99",x"c2",x"49",x"70"),
   438 => (x"fa",x"87",x"c2",x"02"),
   439 => (x"c8",x"49",x"73",x"4c"),
   440 => (x"87",x"ce",x"05",x"99"),
   441 => (x"ff",x"49",x"f5",x"c3"),
   442 => (x"70",x"87",x"eb",x"d5"),
   443 => (x"02",x"99",x"c2",x"49"),
   444 => (x"f8",x"c2",x"87",x"d5"),
   445 => (x"ca",x"02",x"bf",x"f5"),
   446 => (x"88",x"c1",x"48",x"87"),
   447 => (x"58",x"f9",x"f8",x"c2"),
   448 => (x"ff",x"87",x"c2",x"c0"),
   449 => (x"73",x"4d",x"c1",x"4c"),
   450 => (x"05",x"99",x"c4",x"49"),
   451 => (x"f2",x"c3",x"87",x"ce"),
   452 => (x"c1",x"d5",x"ff",x"49"),
   453 => (x"c2",x"49",x"70",x"87"),
   454 => (x"87",x"dc",x"02",x"99"),
   455 => (x"bf",x"f5",x"f8",x"c2"),
   456 => (x"b7",x"c7",x"48",x"7e"),
   457 => (x"cb",x"c0",x"03",x"a8"),
   458 => (x"c1",x"48",x"6e",x"87"),
   459 => (x"f9",x"f8",x"c2",x"80"),
   460 => (x"87",x"c2",x"c0",x"58"),
   461 => (x"4d",x"c1",x"4c",x"fe"),
   462 => (x"ff",x"49",x"fd",x"c3"),
   463 => (x"70",x"87",x"d7",x"d4"),
   464 => (x"02",x"99",x"c2",x"49"),
   465 => (x"c2",x"87",x"d5",x"c0"),
   466 => (x"02",x"bf",x"f5",x"f8"),
   467 => (x"c2",x"87",x"c9",x"c0"),
   468 => (x"c0",x"48",x"f5",x"f8"),
   469 => (x"87",x"c2",x"c0",x"78"),
   470 => (x"4d",x"c1",x"4c",x"fd"),
   471 => (x"ff",x"49",x"fa",x"c3"),
   472 => (x"70",x"87",x"f3",x"d3"),
   473 => (x"02",x"99",x"c2",x"49"),
   474 => (x"c2",x"87",x"d9",x"c0"),
   475 => (x"48",x"bf",x"f5",x"f8"),
   476 => (x"03",x"a8",x"b7",x"c7"),
   477 => (x"c2",x"87",x"c9",x"c0"),
   478 => (x"c7",x"48",x"f5",x"f8"),
   479 => (x"87",x"c2",x"c0",x"78"),
   480 => (x"4d",x"c1",x"4c",x"fc"),
   481 => (x"03",x"ac",x"b7",x"c0"),
   482 => (x"c4",x"87",x"d1",x"c0"),
   483 => (x"d8",x"c1",x"4a",x"66"),
   484 => (x"c0",x"02",x"6a",x"82"),
   485 => (x"4b",x"6a",x"87",x"c6"),
   486 => (x"0f",x"73",x"49",x"74"),
   487 => (x"f0",x"c3",x"1e",x"c0"),
   488 => (x"49",x"da",x"c1",x"1e"),
   489 => (x"c8",x"87",x"ce",x"f7"),
   490 => (x"02",x"98",x"70",x"86"),
   491 => (x"c8",x"87",x"e2",x"c0"),
   492 => (x"f8",x"c2",x"48",x"a6"),
   493 => (x"c8",x"78",x"bf",x"f5"),
   494 => (x"91",x"cb",x"49",x"66"),
   495 => (x"71",x"48",x"66",x"c4"),
   496 => (x"6e",x"7e",x"70",x"80"),
   497 => (x"c8",x"c0",x"02",x"bf"),
   498 => (x"4b",x"bf",x"6e",x"87"),
   499 => (x"73",x"49",x"66",x"c8"),
   500 => (x"02",x"9d",x"75",x"0f"),
   501 => (x"c2",x"87",x"c8",x"c0"),
   502 => (x"49",x"bf",x"f5",x"f8"),
   503 => (x"c2",x"87",x"fa",x"f2"),
   504 => (x"02",x"bf",x"e2",x"e1"),
   505 => (x"49",x"87",x"dd",x"c0"),
   506 => (x"70",x"87",x"c7",x"c2"),
   507 => (x"d3",x"c0",x"02",x"98"),
   508 => (x"f5",x"f8",x"c2",x"87"),
   509 => (x"e0",x"f2",x"49",x"bf"),
   510 => (x"f4",x"49",x"c0",x"87"),
   511 => (x"e1",x"c2",x"87",x"c0"),
   512 => (x"78",x"c0",x"48",x"e2"),
   513 => (x"da",x"f3",x"8e",x"f4"),
   514 => (x"5b",x"5e",x"0e",x"87"),
   515 => (x"1e",x"0e",x"5d",x"5c"),
   516 => (x"f8",x"c2",x"4c",x"71"),
   517 => (x"c1",x"49",x"bf",x"f1"),
   518 => (x"c1",x"4d",x"a1",x"cd"),
   519 => (x"7e",x"69",x"81",x"d1"),
   520 => (x"cf",x"02",x"9c",x"74"),
   521 => (x"4b",x"a5",x"c4",x"87"),
   522 => (x"f8",x"c2",x"7b",x"74"),
   523 => (x"f2",x"49",x"bf",x"f1"),
   524 => (x"7b",x"6e",x"87",x"f9"),
   525 => (x"c4",x"05",x"9c",x"74"),
   526 => (x"c2",x"4b",x"c0",x"87"),
   527 => (x"73",x"4b",x"c1",x"87"),
   528 => (x"87",x"fa",x"f2",x"49"),
   529 => (x"c7",x"02",x"66",x"d4"),
   530 => (x"87",x"da",x"49",x"87"),
   531 => (x"87",x"c2",x"4a",x"70"),
   532 => (x"e1",x"c2",x"4a",x"c0"),
   533 => (x"f2",x"26",x"5a",x"e6"),
   534 => (x"00",x"00",x"87",x"c9"),
   535 => (x"00",x"00",x"00",x"00"),
   536 => (x"00",x"00",x"00",x"00"),
   537 => (x"71",x"1e",x"00",x"00"),
   538 => (x"bf",x"c8",x"ff",x"4a"),
   539 => (x"48",x"a1",x"72",x"49"),
   540 => (x"ff",x"1e",x"4f",x"26"),
   541 => (x"fe",x"89",x"bf",x"c8"),
   542 => (x"c0",x"c0",x"c0",x"c0"),
   543 => (x"c4",x"01",x"a9",x"c0"),
   544 => (x"c2",x"4a",x"c0",x"87"),
   545 => (x"72",x"4a",x"c1",x"87"),
   546 => (x"1e",x"4f",x"26",x"48"),
   547 => (x"bf",x"d9",x"e3",x"c2"),
   548 => (x"c2",x"b9",x"c1",x"49"),
   549 => (x"ff",x"59",x"dd",x"e3"),
   550 => (x"ff",x"c3",x"48",x"d4"),
   551 => (x"48",x"d0",x"ff",x"78"),
   552 => (x"ff",x"78",x"e1",x"c0"),
   553 => (x"78",x"c1",x"48",x"d4"),
   554 => (x"78",x"71",x"31",x"c4"),
   555 => (x"c0",x"48",x"d0",x"ff"),
   556 => (x"4f",x"26",x"78",x"e0"),
   557 => (x"cd",x"e3",x"c2",x"1e"),
   558 => (x"d8",x"f3",x"c2",x"1e"),
   559 => (x"d1",x"fb",x"fd",x"49"),
   560 => (x"70",x"86",x"c4",x"87"),
   561 => (x"87",x"c3",x"02",x"98"),
   562 => (x"26",x"87",x"c0",x"ff"),
   563 => (x"4b",x"35",x"31",x"4f"),
   564 => (x"20",x"20",x"5a",x"48"),
   565 => (x"47",x"46",x"43",x"20"),
   566 => (x"00",x"00",x"00",x"00"),
   567 => (x"5b",x"5e",x"0e",x"00"),
   568 => (x"c2",x"0e",x"5d",x"5c"),
   569 => (x"4a",x"bf",x"e5",x"f8"),
   570 => (x"bf",x"c6",x"e5",x"c2"),
   571 => (x"bc",x"72",x"4c",x"49"),
   572 => (x"c5",x"ff",x"4d",x"71"),
   573 => (x"4b",x"c0",x"87",x"f7"),
   574 => (x"99",x"d0",x"49",x"74"),
   575 => (x"87",x"e7",x"c0",x"02"),
   576 => (x"c8",x"48",x"d0",x"ff"),
   577 => (x"d4",x"ff",x"78",x"e1"),
   578 => (x"75",x"78",x"c5",x"48"),
   579 => (x"02",x"99",x"d0",x"49"),
   580 => (x"f0",x"c3",x"87",x"c3"),
   581 => (x"f4",x"e5",x"c2",x"78"),
   582 => (x"11",x"81",x"73",x"49"),
   583 => (x"08",x"d4",x"ff",x"48"),
   584 => (x"48",x"d0",x"ff",x"78"),
   585 => (x"c1",x"78",x"e0",x"c0"),
   586 => (x"c8",x"83",x"2d",x"2c"),
   587 => (x"c7",x"ff",x"04",x"ab"),
   588 => (x"f0",x"c4",x"ff",x"87"),
   589 => (x"c6",x"e5",x"c2",x"87"),
   590 => (x"e5",x"f8",x"c2",x"48"),
   591 => (x"4d",x"26",x"78",x"bf"),
   592 => (x"4b",x"26",x"4c",x"26"),
   593 => (x"00",x"00",x"4f",x"26"),
   594 => (x"c1",x"1e",x"00",x"00"),
   595 => (x"de",x"48",x"d0",x"e7"),
   596 => (x"dd",x"e5",x"c2",x"50"),
   597 => (x"fa",x"d8",x"fe",x"49"),
   598 => (x"26",x"48",x"c0",x"87"),
   599 => (x"4f",x"54",x"4a",x"4f"),
   600 => (x"55",x"52",x"54",x"55"),
   601 => (x"43",x"52",x"41",x"4e"),
   602 => (x"df",x"f2",x"1e",x"00"),
   603 => (x"87",x"ed",x"fd",x"87"),
   604 => (x"4f",x"26",x"87",x"f8"),
   605 => (x"25",x"26",x"1e",x"16"),
   606 => (x"3e",x"3d",x"36",x"2e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

