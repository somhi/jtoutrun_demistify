
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"fc",x"f8",x"c2",x"87"),
    12 => (x"86",x"c0",x"c5",x"4e"),
    13 => (x"49",x"fc",x"f8",x"c2"),
    14 => (x"48",x"fc",x"e5",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ed",x"e5"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"71",x"1e",x"4f",x"26"),
    53 => (x"49",x"66",x"c4",x"4a"),
    54 => (x"c8",x"88",x"c1",x"48"),
    55 => (x"99",x"71",x"58",x"a6"),
    56 => (x"ff",x"87",x"d6",x"02"),
    57 => (x"ff",x"c3",x"48",x"d4"),
    58 => (x"c4",x"52",x"68",x"78"),
    59 => (x"c1",x"48",x"49",x"66"),
    60 => (x"58",x"a6",x"c8",x"88"),
    61 => (x"ea",x"05",x"99",x"71"),
    62 => (x"1e",x"4f",x"26",x"87"),
    63 => (x"d4",x"ff",x"1e",x"73"),
    64 => (x"7b",x"ff",x"c3",x"4b"),
    65 => (x"ff",x"c3",x"4a",x"6b"),
    66 => (x"c8",x"49",x"6b",x"7b"),
    67 => (x"c3",x"b1",x"72",x"32"),
    68 => (x"4a",x"6b",x"7b",x"ff"),
    69 => (x"b2",x"71",x"31",x"c8"),
    70 => (x"6b",x"7b",x"ff",x"c3"),
    71 => (x"72",x"32",x"c8",x"49"),
    72 => (x"c4",x"48",x"71",x"b1"),
    73 => (x"26",x"4d",x"26",x"87"),
    74 => (x"26",x"4b",x"26",x"4c"),
    75 => (x"5b",x"5e",x"0e",x"4f"),
    76 => (x"71",x"0e",x"5d",x"5c"),
    77 => (x"4c",x"d4",x"ff",x"4a"),
    78 => (x"ff",x"c3",x"49",x"72"),
    79 => (x"c2",x"7c",x"71",x"99"),
    80 => (x"05",x"bf",x"fc",x"e5"),
    81 => (x"66",x"d0",x"87",x"c8"),
    82 => (x"d4",x"30",x"c9",x"48"),
    83 => (x"66",x"d0",x"58",x"a6"),
    84 => (x"c3",x"29",x"d8",x"49"),
    85 => (x"7c",x"71",x"99",x"ff"),
    86 => (x"d0",x"49",x"66",x"d0"),
    87 => (x"99",x"ff",x"c3",x"29"),
    88 => (x"66",x"d0",x"7c",x"71"),
    89 => (x"c3",x"29",x"c8",x"49"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"c3",x"49",x"66",x"d0"),
    92 => (x"7c",x"71",x"99",x"ff"),
    93 => (x"29",x"d0",x"49",x"72"),
    94 => (x"71",x"99",x"ff",x"c3"),
    95 => (x"c9",x"4b",x"6c",x"7c"),
    96 => (x"c3",x"4d",x"ff",x"f0"),
    97 => (x"d0",x"05",x"ab",x"ff"),
    98 => (x"7c",x"ff",x"c3",x"87"),
    99 => (x"8d",x"c1",x"4b",x"6c"),
   100 => (x"c3",x"87",x"c6",x"02"),
   101 => (x"f0",x"02",x"ab",x"ff"),
   102 => (x"fe",x"48",x"73",x"87"),
   103 => (x"c0",x"1e",x"87",x"c7"),
   104 => (x"48",x"d4",x"ff",x"49"),
   105 => (x"c1",x"78",x"ff",x"c3"),
   106 => (x"b7",x"c8",x"c3",x"81"),
   107 => (x"87",x"f1",x"04",x"a9"),
   108 => (x"73",x"1e",x"4f",x"26"),
   109 => (x"c4",x"87",x"e7",x"1e"),
   110 => (x"c0",x"4b",x"df",x"f8"),
   111 => (x"f0",x"ff",x"c0",x"1e"),
   112 => (x"fd",x"49",x"f7",x"c1"),
   113 => (x"86",x"c4",x"87",x"e7"),
   114 => (x"c0",x"05",x"a8",x"c1"),
   115 => (x"d4",x"ff",x"87",x"ea"),
   116 => (x"78",x"ff",x"c3",x"48"),
   117 => (x"c0",x"c0",x"c0",x"c1"),
   118 => (x"c0",x"1e",x"c0",x"c0"),
   119 => (x"e9",x"c1",x"f0",x"e1"),
   120 => (x"87",x"c9",x"fd",x"49"),
   121 => (x"98",x"70",x"86",x"c4"),
   122 => (x"ff",x"87",x"ca",x"05"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"cb",x"48",x"c1",x"78"),
   125 => (x"87",x"e6",x"fe",x"87"),
   126 => (x"fe",x"05",x"8b",x"c1"),
   127 => (x"48",x"c0",x"87",x"fd"),
   128 => (x"1e",x"87",x"e6",x"fc"),
   129 => (x"d4",x"ff",x"1e",x"73"),
   130 => (x"78",x"ff",x"c3",x"48"),
   131 => (x"1e",x"c0",x"4b",x"d3"),
   132 => (x"c1",x"f0",x"ff",x"c0"),
   133 => (x"d4",x"fc",x"49",x"c1"),
   134 => (x"70",x"86",x"c4",x"87"),
   135 => (x"87",x"ca",x"05",x"98"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"48",x"c1",x"78",x"ff"),
   138 => (x"f1",x"fd",x"87",x"cb"),
   139 => (x"05",x"8b",x"c1",x"87"),
   140 => (x"c0",x"87",x"db",x"ff"),
   141 => (x"87",x"f1",x"fb",x"48"),
   142 => (x"5c",x"5b",x"5e",x"0e"),
   143 => (x"4c",x"d4",x"ff",x"0e"),
   144 => (x"c6",x"87",x"db",x"fd"),
   145 => (x"e1",x"c0",x"1e",x"ea"),
   146 => (x"49",x"c8",x"c1",x"f0"),
   147 => (x"c4",x"87",x"de",x"fb"),
   148 => (x"02",x"a8",x"c1",x"86"),
   149 => (x"ea",x"fe",x"87",x"c8"),
   150 => (x"c1",x"48",x"c0",x"87"),
   151 => (x"da",x"fa",x"87",x"e2"),
   152 => (x"cf",x"49",x"70",x"87"),
   153 => (x"c6",x"99",x"ff",x"ff"),
   154 => (x"c8",x"02",x"a9",x"ea"),
   155 => (x"87",x"d3",x"fe",x"87"),
   156 => (x"cb",x"c1",x"48",x"c0"),
   157 => (x"7c",x"ff",x"c3",x"87"),
   158 => (x"fc",x"4b",x"f1",x"c0"),
   159 => (x"98",x"70",x"87",x"f4"),
   160 => (x"87",x"eb",x"c0",x"02"),
   161 => (x"ff",x"c0",x"1e",x"c0"),
   162 => (x"49",x"fa",x"c1",x"f0"),
   163 => (x"c4",x"87",x"de",x"fa"),
   164 => (x"05",x"98",x"70",x"86"),
   165 => (x"ff",x"c3",x"87",x"d9"),
   166 => (x"c3",x"49",x"6c",x"7c"),
   167 => (x"7c",x"7c",x"7c",x"ff"),
   168 => (x"99",x"c0",x"c1",x"7c"),
   169 => (x"c1",x"87",x"c4",x"02"),
   170 => (x"c0",x"87",x"d5",x"48"),
   171 => (x"c2",x"87",x"d1",x"48"),
   172 => (x"87",x"c4",x"05",x"ab"),
   173 => (x"87",x"c8",x"48",x"c0"),
   174 => (x"fe",x"05",x"8b",x"c1"),
   175 => (x"48",x"c0",x"87",x"fd"),
   176 => (x"1e",x"87",x"e4",x"f9"),
   177 => (x"e5",x"c2",x"1e",x"73"),
   178 => (x"78",x"c1",x"48",x"fc"),
   179 => (x"d0",x"ff",x"4b",x"c7"),
   180 => (x"fb",x"78",x"c2",x"48"),
   181 => (x"d0",x"ff",x"87",x"c8"),
   182 => (x"c0",x"78",x"c3",x"48"),
   183 => (x"d0",x"e5",x"c0",x"1e"),
   184 => (x"f9",x"49",x"c0",x"c1"),
   185 => (x"86",x"c4",x"87",x"c7"),
   186 => (x"c1",x"05",x"a8",x"c1"),
   187 => (x"ab",x"c2",x"4b",x"87"),
   188 => (x"c0",x"87",x"c5",x"05"),
   189 => (x"87",x"f9",x"c0",x"48"),
   190 => (x"ff",x"05",x"8b",x"c1"),
   191 => (x"f7",x"fc",x"87",x"d0"),
   192 => (x"c0",x"e6",x"c2",x"87"),
   193 => (x"05",x"98",x"70",x"58"),
   194 => (x"1e",x"c1",x"87",x"cd"),
   195 => (x"c1",x"f0",x"ff",x"c0"),
   196 => (x"d8",x"f8",x"49",x"d0"),
   197 => (x"ff",x"86",x"c4",x"87"),
   198 => (x"ff",x"c3",x"48",x"d4"),
   199 => (x"87",x"fc",x"c2",x"78"),
   200 => (x"58",x"c4",x"e6",x"c2"),
   201 => (x"c2",x"48",x"d0",x"ff"),
   202 => (x"48",x"d4",x"ff",x"78"),
   203 => (x"c1",x"78",x"ff",x"c3"),
   204 => (x"87",x"f5",x"f7",x"48"),
   205 => (x"5c",x"5b",x"5e",x"0e"),
   206 => (x"4b",x"71",x"0e",x"5d"),
   207 => (x"ee",x"c5",x"4c",x"c0"),
   208 => (x"ff",x"4a",x"df",x"cd"),
   209 => (x"ff",x"c3",x"48",x"d4"),
   210 => (x"c3",x"49",x"68",x"78"),
   211 => (x"c0",x"05",x"a9",x"fe"),
   212 => (x"4d",x"70",x"87",x"fd"),
   213 => (x"cc",x"02",x"9b",x"73"),
   214 => (x"1e",x"66",x"d0",x"87"),
   215 => (x"f1",x"f5",x"49",x"73"),
   216 => (x"d6",x"86",x"c4",x"87"),
   217 => (x"48",x"d0",x"ff",x"87"),
   218 => (x"c3",x"78",x"d1",x"c4"),
   219 => (x"66",x"d0",x"7d",x"ff"),
   220 => (x"d4",x"88",x"c1",x"48"),
   221 => (x"98",x"70",x"58",x"a6"),
   222 => (x"ff",x"87",x"f0",x"05"),
   223 => (x"ff",x"c3",x"48",x"d4"),
   224 => (x"9b",x"73",x"78",x"78"),
   225 => (x"ff",x"87",x"c5",x"05"),
   226 => (x"78",x"d0",x"48",x"d0"),
   227 => (x"c1",x"4c",x"4a",x"c1"),
   228 => (x"ee",x"fe",x"05",x"8a"),
   229 => (x"f6",x"48",x"74",x"87"),
   230 => (x"73",x"1e",x"87",x"cb"),
   231 => (x"c0",x"4a",x"71",x"1e"),
   232 => (x"48",x"d4",x"ff",x"4b"),
   233 => (x"ff",x"78",x"ff",x"c3"),
   234 => (x"c3",x"c4",x"48",x"d0"),
   235 => (x"48",x"d4",x"ff",x"78"),
   236 => (x"72",x"78",x"ff",x"c3"),
   237 => (x"f0",x"ff",x"c0",x"1e"),
   238 => (x"f5",x"49",x"d1",x"c1"),
   239 => (x"86",x"c4",x"87",x"ef"),
   240 => (x"d2",x"05",x"98",x"70"),
   241 => (x"1e",x"c0",x"c8",x"87"),
   242 => (x"fd",x"49",x"66",x"cc"),
   243 => (x"86",x"c4",x"87",x"e6"),
   244 => (x"d0",x"ff",x"4b",x"70"),
   245 => (x"73",x"78",x"c2",x"48"),
   246 => (x"87",x"cd",x"f5",x"48"),
   247 => (x"5c",x"5b",x"5e",x"0e"),
   248 => (x"1e",x"c0",x"0e",x"5d"),
   249 => (x"c1",x"f0",x"ff",x"c0"),
   250 => (x"c0",x"f5",x"49",x"c9"),
   251 => (x"c2",x"1e",x"d2",x"87"),
   252 => (x"fc",x"49",x"c4",x"e6"),
   253 => (x"86",x"c8",x"87",x"fe"),
   254 => (x"84",x"c1",x"4c",x"c0"),
   255 => (x"04",x"ac",x"b7",x"d2"),
   256 => (x"e6",x"c2",x"87",x"f8"),
   257 => (x"49",x"bf",x"97",x"c4"),
   258 => (x"c1",x"99",x"c0",x"c3"),
   259 => (x"c0",x"05",x"a9",x"c0"),
   260 => (x"e6",x"c2",x"87",x"e7"),
   261 => (x"49",x"bf",x"97",x"cb"),
   262 => (x"e6",x"c2",x"31",x"d0"),
   263 => (x"4a",x"bf",x"97",x"cc"),
   264 => (x"b1",x"72",x"32",x"c8"),
   265 => (x"97",x"cd",x"e6",x"c2"),
   266 => (x"71",x"b1",x"4a",x"bf"),
   267 => (x"ff",x"ff",x"cf",x"4c"),
   268 => (x"84",x"c1",x"9c",x"ff"),
   269 => (x"e7",x"c1",x"34",x"ca"),
   270 => (x"cd",x"e6",x"c2",x"87"),
   271 => (x"c1",x"49",x"bf",x"97"),
   272 => (x"c2",x"99",x"c6",x"31"),
   273 => (x"bf",x"97",x"ce",x"e6"),
   274 => (x"2a",x"b7",x"c7",x"4a"),
   275 => (x"e6",x"c2",x"b1",x"72"),
   276 => (x"4a",x"bf",x"97",x"c9"),
   277 => (x"c2",x"9d",x"cf",x"4d"),
   278 => (x"bf",x"97",x"ca",x"e6"),
   279 => (x"ca",x"9a",x"c3",x"4a"),
   280 => (x"cb",x"e6",x"c2",x"32"),
   281 => (x"c2",x"4b",x"bf",x"97"),
   282 => (x"c2",x"b2",x"73",x"33"),
   283 => (x"bf",x"97",x"cc",x"e6"),
   284 => (x"9b",x"c0",x"c3",x"4b"),
   285 => (x"73",x"2b",x"b7",x"c6"),
   286 => (x"c1",x"81",x"c2",x"b2"),
   287 => (x"70",x"30",x"71",x"48"),
   288 => (x"75",x"48",x"c1",x"49"),
   289 => (x"72",x"4d",x"70",x"30"),
   290 => (x"71",x"84",x"c1",x"4c"),
   291 => (x"b7",x"c0",x"c8",x"94"),
   292 => (x"87",x"cc",x"06",x"ad"),
   293 => (x"2d",x"b7",x"34",x"c1"),
   294 => (x"ad",x"b7",x"c0",x"c8"),
   295 => (x"87",x"f4",x"ff",x"01"),
   296 => (x"c0",x"f2",x"48",x"74"),
   297 => (x"5b",x"5e",x"0e",x"87"),
   298 => (x"f8",x"0e",x"5d",x"5c"),
   299 => (x"ea",x"ee",x"c2",x"86"),
   300 => (x"c2",x"78",x"c0",x"48"),
   301 => (x"c0",x"1e",x"e2",x"e6"),
   302 => (x"87",x"de",x"fb",x"49"),
   303 => (x"98",x"70",x"86",x"c4"),
   304 => (x"c0",x"87",x"c5",x"05"),
   305 => (x"87",x"ce",x"c9",x"48"),
   306 => (x"7e",x"c1",x"4d",x"c0"),
   307 => (x"bf",x"e1",x"f5",x"c0"),
   308 => (x"d8",x"e7",x"c2",x"49"),
   309 => (x"4b",x"c8",x"71",x"4a"),
   310 => (x"70",x"87",x"cf",x"ee"),
   311 => (x"87",x"c2",x"05",x"98"),
   312 => (x"f5",x"c0",x"7e",x"c0"),
   313 => (x"c2",x"49",x"bf",x"dd"),
   314 => (x"71",x"4a",x"f4",x"e7"),
   315 => (x"f9",x"ed",x"4b",x"c8"),
   316 => (x"05",x"98",x"70",x"87"),
   317 => (x"7e",x"c0",x"87",x"c2"),
   318 => (x"fd",x"c0",x"02",x"6e"),
   319 => (x"e8",x"ed",x"c2",x"87"),
   320 => (x"ee",x"c2",x"4d",x"bf"),
   321 => (x"7e",x"bf",x"9f",x"e0"),
   322 => (x"ea",x"d6",x"c5",x"48"),
   323 => (x"87",x"c7",x"05",x"a8"),
   324 => (x"bf",x"e8",x"ed",x"c2"),
   325 => (x"6e",x"87",x"ce",x"4d"),
   326 => (x"d5",x"e9",x"ca",x"48"),
   327 => (x"87",x"c5",x"02",x"a8"),
   328 => (x"f1",x"c7",x"48",x"c0"),
   329 => (x"e2",x"e6",x"c2",x"87"),
   330 => (x"f9",x"49",x"75",x"1e"),
   331 => (x"86",x"c4",x"87",x"ec"),
   332 => (x"c5",x"05",x"98",x"70"),
   333 => (x"c7",x"48",x"c0",x"87"),
   334 => (x"f5",x"c0",x"87",x"dc"),
   335 => (x"c2",x"49",x"bf",x"dd"),
   336 => (x"71",x"4a",x"f4",x"e7"),
   337 => (x"e1",x"ec",x"4b",x"c8"),
   338 => (x"05",x"98",x"70",x"87"),
   339 => (x"ee",x"c2",x"87",x"c8"),
   340 => (x"78",x"c1",x"48",x"ea"),
   341 => (x"f5",x"c0",x"87",x"da"),
   342 => (x"c2",x"49",x"bf",x"e1"),
   343 => (x"71",x"4a",x"d8",x"e7"),
   344 => (x"c5",x"ec",x"4b",x"c8"),
   345 => (x"02",x"98",x"70",x"87"),
   346 => (x"c0",x"87",x"c5",x"c0"),
   347 => (x"87",x"e6",x"c6",x"48"),
   348 => (x"97",x"e0",x"ee",x"c2"),
   349 => (x"d5",x"c1",x"49",x"bf"),
   350 => (x"cd",x"c0",x"05",x"a9"),
   351 => (x"e1",x"ee",x"c2",x"87"),
   352 => (x"c2",x"49",x"bf",x"97"),
   353 => (x"c0",x"02",x"a9",x"ea"),
   354 => (x"48",x"c0",x"87",x"c5"),
   355 => (x"c2",x"87",x"c7",x"c6"),
   356 => (x"bf",x"97",x"e2",x"e6"),
   357 => (x"e9",x"c3",x"48",x"7e"),
   358 => (x"ce",x"c0",x"02",x"a8"),
   359 => (x"c3",x"48",x"6e",x"87"),
   360 => (x"c0",x"02",x"a8",x"eb"),
   361 => (x"48",x"c0",x"87",x"c5"),
   362 => (x"c2",x"87",x"eb",x"c5"),
   363 => (x"bf",x"97",x"ed",x"e6"),
   364 => (x"c0",x"05",x"99",x"49"),
   365 => (x"e6",x"c2",x"87",x"cc"),
   366 => (x"49",x"bf",x"97",x"ee"),
   367 => (x"c0",x"02",x"a9",x"c2"),
   368 => (x"48",x"c0",x"87",x"c5"),
   369 => (x"c2",x"87",x"cf",x"c5"),
   370 => (x"bf",x"97",x"ef",x"e6"),
   371 => (x"e6",x"ee",x"c2",x"48"),
   372 => (x"48",x"4c",x"70",x"58"),
   373 => (x"ee",x"c2",x"88",x"c1"),
   374 => (x"e6",x"c2",x"58",x"ea"),
   375 => (x"49",x"bf",x"97",x"f0"),
   376 => (x"e6",x"c2",x"81",x"75"),
   377 => (x"4a",x"bf",x"97",x"f1"),
   378 => (x"a1",x"72",x"32",x"c8"),
   379 => (x"f7",x"f2",x"c2",x"7e"),
   380 => (x"c2",x"78",x"6e",x"48"),
   381 => (x"bf",x"97",x"f2",x"e6"),
   382 => (x"58",x"a6",x"c8",x"48"),
   383 => (x"bf",x"ea",x"ee",x"c2"),
   384 => (x"87",x"d4",x"c2",x"02"),
   385 => (x"bf",x"dd",x"f5",x"c0"),
   386 => (x"f4",x"e7",x"c2",x"49"),
   387 => (x"4b",x"c8",x"71",x"4a"),
   388 => (x"70",x"87",x"d7",x"e9"),
   389 => (x"c5",x"c0",x"02",x"98"),
   390 => (x"c3",x"48",x"c0",x"87"),
   391 => (x"ee",x"c2",x"87",x"f8"),
   392 => (x"c2",x"4c",x"bf",x"e2"),
   393 => (x"c2",x"5c",x"cb",x"f3"),
   394 => (x"bf",x"97",x"c7",x"e7"),
   395 => (x"c2",x"31",x"c8",x"49"),
   396 => (x"bf",x"97",x"c6",x"e7"),
   397 => (x"c2",x"49",x"a1",x"4a"),
   398 => (x"bf",x"97",x"c8",x"e7"),
   399 => (x"72",x"32",x"d0",x"4a"),
   400 => (x"e7",x"c2",x"49",x"a1"),
   401 => (x"4a",x"bf",x"97",x"c9"),
   402 => (x"a1",x"72",x"32",x"d8"),
   403 => (x"91",x"66",x"c4",x"49"),
   404 => (x"bf",x"f7",x"f2",x"c2"),
   405 => (x"ff",x"f2",x"c2",x"81"),
   406 => (x"cf",x"e7",x"c2",x"59"),
   407 => (x"c8",x"4a",x"bf",x"97"),
   408 => (x"ce",x"e7",x"c2",x"32"),
   409 => (x"a2",x"4b",x"bf",x"97"),
   410 => (x"d0",x"e7",x"c2",x"4a"),
   411 => (x"d0",x"4b",x"bf",x"97"),
   412 => (x"4a",x"a2",x"73",x"33"),
   413 => (x"97",x"d1",x"e7",x"c2"),
   414 => (x"9b",x"cf",x"4b",x"bf"),
   415 => (x"a2",x"73",x"33",x"d8"),
   416 => (x"c3",x"f3",x"c2",x"4a"),
   417 => (x"ff",x"f2",x"c2",x"5a"),
   418 => (x"8a",x"c2",x"4a",x"bf"),
   419 => (x"f3",x"c2",x"92",x"74"),
   420 => (x"a1",x"72",x"48",x"c3"),
   421 => (x"87",x"ca",x"c1",x"78"),
   422 => (x"97",x"f4",x"e6",x"c2"),
   423 => (x"31",x"c8",x"49",x"bf"),
   424 => (x"97",x"f3",x"e6",x"c2"),
   425 => (x"49",x"a1",x"4a",x"bf"),
   426 => (x"59",x"f2",x"ee",x"c2"),
   427 => (x"bf",x"ee",x"ee",x"c2"),
   428 => (x"c7",x"31",x"c5",x"49"),
   429 => (x"29",x"c9",x"81",x"ff"),
   430 => (x"59",x"cb",x"f3",x"c2"),
   431 => (x"97",x"f9",x"e6",x"c2"),
   432 => (x"32",x"c8",x"4a",x"bf"),
   433 => (x"97",x"f8",x"e6",x"c2"),
   434 => (x"4a",x"a2",x"4b",x"bf"),
   435 => (x"6e",x"92",x"66",x"c4"),
   436 => (x"c7",x"f3",x"c2",x"82"),
   437 => (x"ff",x"f2",x"c2",x"5a"),
   438 => (x"c2",x"78",x"c0",x"48"),
   439 => (x"72",x"48",x"fb",x"f2"),
   440 => (x"f3",x"c2",x"78",x"a1"),
   441 => (x"f2",x"c2",x"48",x"cb"),
   442 => (x"c2",x"78",x"bf",x"ff"),
   443 => (x"c2",x"48",x"cf",x"f3"),
   444 => (x"78",x"bf",x"c3",x"f3"),
   445 => (x"bf",x"ea",x"ee",x"c2"),
   446 => (x"87",x"c9",x"c0",x"02"),
   447 => (x"30",x"c4",x"48",x"74"),
   448 => (x"c9",x"c0",x"7e",x"70"),
   449 => (x"c7",x"f3",x"c2",x"87"),
   450 => (x"30",x"c4",x"48",x"bf"),
   451 => (x"ee",x"c2",x"7e",x"70"),
   452 => (x"78",x"6e",x"48",x"ee"),
   453 => (x"8e",x"f8",x"48",x"c1"),
   454 => (x"4c",x"26",x"4d",x"26"),
   455 => (x"4f",x"26",x"4b",x"26"),
   456 => (x"5c",x"5b",x"5e",x"0e"),
   457 => (x"4a",x"71",x"0e",x"5d"),
   458 => (x"bf",x"ea",x"ee",x"c2"),
   459 => (x"72",x"87",x"cb",x"02"),
   460 => (x"72",x"2b",x"c7",x"4b"),
   461 => (x"9c",x"ff",x"c1",x"4c"),
   462 => (x"4b",x"72",x"87",x"c9"),
   463 => (x"4c",x"72",x"2b",x"c8"),
   464 => (x"c2",x"9c",x"ff",x"c3"),
   465 => (x"83",x"bf",x"f7",x"f2"),
   466 => (x"bf",x"d9",x"f5",x"c0"),
   467 => (x"87",x"d9",x"02",x"ab"),
   468 => (x"5b",x"dd",x"f5",x"c0"),
   469 => (x"1e",x"e2",x"e6",x"c2"),
   470 => (x"fd",x"f0",x"49",x"73"),
   471 => (x"70",x"86",x"c4",x"87"),
   472 => (x"87",x"c5",x"05",x"98"),
   473 => (x"e6",x"c0",x"48",x"c0"),
   474 => (x"ea",x"ee",x"c2",x"87"),
   475 => (x"87",x"d2",x"02",x"bf"),
   476 => (x"91",x"c4",x"49",x"74"),
   477 => (x"81",x"e2",x"e6",x"c2"),
   478 => (x"ff",x"cf",x"4d",x"69"),
   479 => (x"9d",x"ff",x"ff",x"ff"),
   480 => (x"49",x"74",x"87",x"cb"),
   481 => (x"e6",x"c2",x"91",x"c2"),
   482 => (x"69",x"9f",x"81",x"e2"),
   483 => (x"fe",x"48",x"75",x"4d"),
   484 => (x"5e",x"0e",x"87",x"c6"),
   485 => (x"0e",x"5d",x"5c",x"5b"),
   486 => (x"4c",x"71",x"86",x"f8"),
   487 => (x"87",x"c5",x"05",x"9c"),
   488 => (x"c1",x"c3",x"48",x"c0"),
   489 => (x"7e",x"a4",x"c8",x"87"),
   490 => (x"78",x"c0",x"48",x"6e"),
   491 => (x"c7",x"02",x"66",x"d8"),
   492 => (x"97",x"66",x"d8",x"87"),
   493 => (x"87",x"c5",x"05",x"bf"),
   494 => (x"e9",x"c2",x"48",x"c0"),
   495 => (x"c1",x"1e",x"c0",x"87"),
   496 => (x"87",x"f9",x"ce",x"49"),
   497 => (x"4d",x"70",x"86",x"c4"),
   498 => (x"c2",x"c1",x"02",x"9d"),
   499 => (x"f2",x"ee",x"c2",x"87"),
   500 => (x"49",x"66",x"d8",x"4a"),
   501 => (x"70",x"87",x"f8",x"e1"),
   502 => (x"f2",x"c0",x"02",x"98"),
   503 => (x"d8",x"4a",x"75",x"87"),
   504 => (x"4b",x"cb",x"49",x"66"),
   505 => (x"70",x"87",x"dd",x"e2"),
   506 => (x"e2",x"c0",x"02",x"98"),
   507 => (x"75",x"1e",x"c0",x"87"),
   508 => (x"87",x"c7",x"02",x"9d"),
   509 => (x"c0",x"48",x"a6",x"c8"),
   510 => (x"c8",x"87",x"c5",x"78"),
   511 => (x"78",x"c1",x"48",x"a6"),
   512 => (x"cd",x"49",x"66",x"c8"),
   513 => (x"86",x"c4",x"87",x"f7"),
   514 => (x"05",x"9d",x"4d",x"70"),
   515 => (x"75",x"87",x"fe",x"fe"),
   516 => (x"cf",x"c1",x"02",x"9d"),
   517 => (x"49",x"a5",x"dc",x"87"),
   518 => (x"78",x"69",x"48",x"6e"),
   519 => (x"c4",x"49",x"a5",x"da"),
   520 => (x"a4",x"c4",x"48",x"a6"),
   521 => (x"48",x"69",x"9f",x"78"),
   522 => (x"78",x"08",x"66",x"c4"),
   523 => (x"bf",x"ea",x"ee",x"c2"),
   524 => (x"d4",x"87",x"d2",x"02"),
   525 => (x"69",x"9f",x"49",x"a5"),
   526 => (x"ff",x"ff",x"c0",x"49"),
   527 => (x"d0",x"48",x"71",x"99"),
   528 => (x"c2",x"7e",x"70",x"30"),
   529 => (x"6e",x"7e",x"c0",x"87"),
   530 => (x"66",x"c4",x"48",x"49"),
   531 => (x"66",x"c4",x"80",x"bf"),
   532 => (x"7c",x"c0",x"78",x"08"),
   533 => (x"c4",x"49",x"a4",x"cc"),
   534 => (x"d0",x"79",x"bf",x"66"),
   535 => (x"79",x"c0",x"49",x"a4"),
   536 => (x"87",x"c2",x"48",x"c1"),
   537 => (x"8e",x"f8",x"48",x"c0"),
   538 => (x"0e",x"87",x"ed",x"fa"),
   539 => (x"5d",x"5c",x"5b",x"5e"),
   540 => (x"9c",x"4c",x"71",x"0e"),
   541 => (x"87",x"ca",x"c1",x"02"),
   542 => (x"69",x"49",x"a4",x"c8"),
   543 => (x"87",x"c2",x"c1",x"02"),
   544 => (x"6c",x"4a",x"66",x"d0"),
   545 => (x"a6",x"d4",x"82",x"49"),
   546 => (x"4d",x"66",x"d0",x"5a"),
   547 => (x"e6",x"ee",x"c2",x"b9"),
   548 => (x"ba",x"ff",x"4a",x"bf"),
   549 => (x"99",x"71",x"99",x"72"),
   550 => (x"87",x"e4",x"c0",x"02"),
   551 => (x"6b",x"4b",x"a4",x"c4"),
   552 => (x"87",x"fc",x"f9",x"49"),
   553 => (x"ee",x"c2",x"7b",x"70"),
   554 => (x"6c",x"49",x"bf",x"e2"),
   555 => (x"75",x"7c",x"71",x"81"),
   556 => (x"e6",x"ee",x"c2",x"b9"),
   557 => (x"ba",x"ff",x"4a",x"bf"),
   558 => (x"99",x"71",x"99",x"72"),
   559 => (x"87",x"dc",x"ff",x"05"),
   560 => (x"d3",x"f9",x"7c",x"75"),
   561 => (x"1e",x"73",x"1e",x"87"),
   562 => (x"02",x"9b",x"4b",x"71"),
   563 => (x"a3",x"c8",x"87",x"c7"),
   564 => (x"c5",x"05",x"69",x"49"),
   565 => (x"c0",x"48",x"c0",x"87"),
   566 => (x"f2",x"c2",x"87",x"f7"),
   567 => (x"c4",x"4a",x"bf",x"fb"),
   568 => (x"49",x"69",x"49",x"a3"),
   569 => (x"ee",x"c2",x"89",x"c2"),
   570 => (x"71",x"91",x"bf",x"e2"),
   571 => (x"ee",x"c2",x"4a",x"a2"),
   572 => (x"6b",x"49",x"bf",x"e6"),
   573 => (x"4a",x"a2",x"71",x"99"),
   574 => (x"5a",x"dd",x"f5",x"c0"),
   575 => (x"72",x"1e",x"66",x"c8"),
   576 => (x"87",x"d6",x"ea",x"49"),
   577 => (x"98",x"70",x"86",x"c4"),
   578 => (x"c0",x"87",x"c4",x"05"),
   579 => (x"c1",x"87",x"c2",x"48"),
   580 => (x"87",x"c8",x"f8",x"48"),
   581 => (x"5c",x"5b",x"5e",x"0e"),
   582 => (x"71",x"1e",x"0e",x"5d"),
   583 => (x"4c",x"66",x"d4",x"4b"),
   584 => (x"9b",x"73",x"2c",x"c9"),
   585 => (x"87",x"cf",x"c1",x"02"),
   586 => (x"69",x"49",x"a3",x"c8"),
   587 => (x"87",x"c7",x"c1",x"02"),
   588 => (x"d4",x"4d",x"a3",x"d0"),
   589 => (x"ee",x"c2",x"7d",x"66"),
   590 => (x"ff",x"49",x"bf",x"e6"),
   591 => (x"99",x"4a",x"6b",x"b9"),
   592 => (x"03",x"ac",x"71",x"7e"),
   593 => (x"7b",x"c0",x"87",x"cd"),
   594 => (x"4a",x"a3",x"cc",x"7d"),
   595 => (x"6a",x"49",x"a3",x"c4"),
   596 => (x"72",x"87",x"c2",x"79"),
   597 => (x"02",x"9c",x"74",x"8c"),
   598 => (x"1e",x"49",x"87",x"dd"),
   599 => (x"ca",x"fc",x"49",x"73"),
   600 => (x"d4",x"86",x"c4",x"87"),
   601 => (x"ff",x"c7",x"49",x"66"),
   602 => (x"87",x"cb",x"02",x"99"),
   603 => (x"1e",x"e2",x"e6",x"c2"),
   604 => (x"d0",x"fd",x"49",x"73"),
   605 => (x"26",x"86",x"c4",x"87"),
   606 => (x"0e",x"87",x"dd",x"f6"),
   607 => (x"5d",x"5c",x"5b",x"5e"),
   608 => (x"d0",x"86",x"f0",x"0e"),
   609 => (x"e4",x"c0",x"59",x"a6"),
   610 => (x"66",x"cc",x"4b",x"66"),
   611 => (x"48",x"87",x"ca",x"02"),
   612 => (x"7e",x"70",x"80",x"c8"),
   613 => (x"c5",x"05",x"bf",x"6e"),
   614 => (x"c3",x"48",x"c0",x"87"),
   615 => (x"66",x"cc",x"87",x"ec"),
   616 => (x"73",x"84",x"d0",x"4c"),
   617 => (x"48",x"a6",x"c4",x"49"),
   618 => (x"66",x"c4",x"78",x"6c"),
   619 => (x"6e",x"80",x"c4",x"81"),
   620 => (x"66",x"c8",x"78",x"bf"),
   621 => (x"87",x"c6",x"06",x"a9"),
   622 => (x"89",x"66",x"c4",x"49"),
   623 => (x"b7",x"c0",x"4b",x"71"),
   624 => (x"87",x"c4",x"01",x"ab"),
   625 => (x"87",x"c2",x"c3",x"48"),
   626 => (x"c7",x"48",x"66",x"c4"),
   627 => (x"7e",x"70",x"98",x"ff"),
   628 => (x"c9",x"c1",x"02",x"6e"),
   629 => (x"49",x"c0",x"c8",x"87"),
   630 => (x"4a",x"71",x"89",x"6e"),
   631 => (x"4d",x"e2",x"e6",x"c2"),
   632 => (x"b7",x"73",x"85",x"6e"),
   633 => (x"87",x"c1",x"06",x"aa"),
   634 => (x"48",x"49",x"72",x"4a"),
   635 => (x"70",x"80",x"66",x"c4"),
   636 => (x"49",x"8b",x"72",x"7c"),
   637 => (x"99",x"71",x"8a",x"c1"),
   638 => (x"c0",x"87",x"d9",x"02"),
   639 => (x"15",x"48",x"66",x"e0"),
   640 => (x"66",x"e0",x"c0",x"50"),
   641 => (x"c0",x"80",x"c1",x"48"),
   642 => (x"72",x"58",x"a6",x"e4"),
   643 => (x"71",x"8a",x"c1",x"49"),
   644 => (x"87",x"e7",x"05",x"99"),
   645 => (x"66",x"d0",x"1e",x"c1"),
   646 => (x"87",x"cf",x"f9",x"49"),
   647 => (x"b7",x"c0",x"86",x"c4"),
   648 => (x"e3",x"c1",x"06",x"ab"),
   649 => (x"66",x"e0",x"c0",x"87"),
   650 => (x"b7",x"ff",x"c7",x"4d"),
   651 => (x"e2",x"c0",x"06",x"ab"),
   652 => (x"d0",x"1e",x"75",x"87"),
   653 => (x"cc",x"fa",x"49",x"66"),
   654 => (x"85",x"c0",x"c8",x"87"),
   655 => (x"c0",x"c8",x"48",x"6c"),
   656 => (x"c8",x"7c",x"70",x"80"),
   657 => (x"1e",x"c1",x"8b",x"c0"),
   658 => (x"f8",x"49",x"66",x"d4"),
   659 => (x"86",x"c8",x"87",x"dd"),
   660 => (x"c2",x"87",x"ee",x"c0"),
   661 => (x"d0",x"1e",x"e2",x"e6"),
   662 => (x"e8",x"f9",x"49",x"66"),
   663 => (x"c2",x"86",x"c4",x"87"),
   664 => (x"73",x"4a",x"e2",x"e6"),
   665 => (x"80",x"6c",x"48",x"49"),
   666 => (x"49",x"73",x"7c",x"70"),
   667 => (x"99",x"71",x"8b",x"c1"),
   668 => (x"12",x"87",x"ce",x"02"),
   669 => (x"85",x"c1",x"7d",x"97"),
   670 => (x"8b",x"c1",x"49",x"73"),
   671 => (x"f2",x"05",x"99",x"71"),
   672 => (x"ab",x"b7",x"c0",x"87"),
   673 => (x"87",x"e1",x"fe",x"01"),
   674 => (x"8e",x"f0",x"48",x"c1"),
   675 => (x"0e",x"87",x"c9",x"f2"),
   676 => (x"5d",x"5c",x"5b",x"5e"),
   677 => (x"9b",x"4b",x"71",x"0e"),
   678 => (x"c8",x"87",x"c7",x"02"),
   679 => (x"05",x"6d",x"4d",x"a3"),
   680 => (x"48",x"ff",x"87",x"c5"),
   681 => (x"d0",x"87",x"fd",x"c0"),
   682 => (x"49",x"6c",x"4c",x"a3"),
   683 => (x"05",x"99",x"ff",x"c7"),
   684 => (x"02",x"6c",x"87",x"d8"),
   685 => (x"1e",x"c1",x"87",x"c9"),
   686 => (x"ee",x"f6",x"49",x"73"),
   687 => (x"c2",x"86",x"c4",x"87"),
   688 => (x"73",x"1e",x"e2",x"e6"),
   689 => (x"87",x"fd",x"f7",x"49"),
   690 => (x"4a",x"6c",x"86",x"c4"),
   691 => (x"c4",x"04",x"aa",x"6d"),
   692 => (x"cf",x"48",x"ff",x"87"),
   693 => (x"7c",x"a2",x"c1",x"87"),
   694 => (x"ff",x"c7",x"49",x"72"),
   695 => (x"e2",x"e6",x"c2",x"99"),
   696 => (x"48",x"69",x"97",x"81"),
   697 => (x"1e",x"87",x"f1",x"f0"),
   698 => (x"4b",x"71",x"1e",x"73"),
   699 => (x"e4",x"c0",x"02",x"9b"),
   700 => (x"cf",x"f3",x"c2",x"87"),
   701 => (x"c2",x"4a",x"73",x"5b"),
   702 => (x"e2",x"ee",x"c2",x"8a"),
   703 => (x"c2",x"92",x"49",x"bf"),
   704 => (x"48",x"bf",x"fb",x"f2"),
   705 => (x"f3",x"c2",x"80",x"72"),
   706 => (x"48",x"71",x"58",x"d3"),
   707 => (x"ee",x"c2",x"30",x"c4"),
   708 => (x"ed",x"c0",x"58",x"f2"),
   709 => (x"cb",x"f3",x"c2",x"87"),
   710 => (x"ff",x"f2",x"c2",x"48"),
   711 => (x"f3",x"c2",x"78",x"bf"),
   712 => (x"f3",x"c2",x"48",x"cf"),
   713 => (x"c2",x"78",x"bf",x"c3"),
   714 => (x"02",x"bf",x"ea",x"ee"),
   715 => (x"ee",x"c2",x"87",x"c9"),
   716 => (x"c4",x"49",x"bf",x"e2"),
   717 => (x"c2",x"87",x"c7",x"31"),
   718 => (x"49",x"bf",x"c7",x"f3"),
   719 => (x"ee",x"c2",x"31",x"c4"),
   720 => (x"d7",x"ef",x"59",x"f2"),
   721 => (x"5b",x"5e",x"0e",x"87"),
   722 => (x"4a",x"71",x"0e",x"5c"),
   723 => (x"9a",x"72",x"4b",x"c0"),
   724 => (x"87",x"e1",x"c0",x"02"),
   725 => (x"9f",x"49",x"a2",x"da"),
   726 => (x"ee",x"c2",x"4b",x"69"),
   727 => (x"cf",x"02",x"bf",x"ea"),
   728 => (x"49",x"a2",x"d4",x"87"),
   729 => (x"4c",x"49",x"69",x"9f"),
   730 => (x"9c",x"ff",x"ff",x"c0"),
   731 => (x"87",x"c2",x"34",x"d0"),
   732 => (x"49",x"74",x"4c",x"c0"),
   733 => (x"fd",x"49",x"73",x"b3"),
   734 => (x"dd",x"ee",x"87",x"ed"),
   735 => (x"5b",x"5e",x"0e",x"87"),
   736 => (x"f4",x"0e",x"5d",x"5c"),
   737 => (x"c0",x"4a",x"71",x"86"),
   738 => (x"02",x"9a",x"72",x"7e"),
   739 => (x"e6",x"c2",x"87",x"d8"),
   740 => (x"78",x"c0",x"48",x"de"),
   741 => (x"48",x"d6",x"e6",x"c2"),
   742 => (x"bf",x"cf",x"f3",x"c2"),
   743 => (x"da",x"e6",x"c2",x"78"),
   744 => (x"cb",x"f3",x"c2",x"48"),
   745 => (x"ee",x"c2",x"78",x"bf"),
   746 => (x"50",x"c0",x"48",x"ff"),
   747 => (x"bf",x"ee",x"ee",x"c2"),
   748 => (x"de",x"e6",x"c2",x"49"),
   749 => (x"aa",x"71",x"4a",x"bf"),
   750 => (x"87",x"ca",x"c4",x"03"),
   751 => (x"99",x"cf",x"49",x"72"),
   752 => (x"87",x"ea",x"c0",x"05"),
   753 => (x"48",x"d9",x"f5",x"c0"),
   754 => (x"bf",x"d6",x"e6",x"c2"),
   755 => (x"e2",x"e6",x"c2",x"78"),
   756 => (x"d6",x"e6",x"c2",x"1e"),
   757 => (x"e6",x"c2",x"49",x"bf"),
   758 => (x"a1",x"c1",x"48",x"d6"),
   759 => (x"de",x"ff",x"71",x"78"),
   760 => (x"86",x"c4",x"87",x"f8"),
   761 => (x"48",x"d5",x"f5",x"c0"),
   762 => (x"78",x"e2",x"e6",x"c2"),
   763 => (x"f5",x"c0",x"87",x"cc"),
   764 => (x"c0",x"48",x"bf",x"d5"),
   765 => (x"f5",x"c0",x"80",x"e0"),
   766 => (x"e6",x"c2",x"58",x"d9"),
   767 => (x"c1",x"48",x"bf",x"de"),
   768 => (x"e2",x"e6",x"c2",x"80"),
   769 => (x"0d",x"55",x"27",x"58"),
   770 => (x"97",x"bf",x"00",x"00"),
   771 => (x"02",x"9d",x"4d",x"bf"),
   772 => (x"c3",x"87",x"e3",x"c2"),
   773 => (x"c2",x"02",x"ad",x"e5"),
   774 => (x"f5",x"c0",x"87",x"dc"),
   775 => (x"cb",x"4b",x"bf",x"d5"),
   776 => (x"4c",x"11",x"49",x"a3"),
   777 => (x"c1",x"05",x"ac",x"cf"),
   778 => (x"49",x"75",x"87",x"d2"),
   779 => (x"89",x"c1",x"99",x"df"),
   780 => (x"ee",x"c2",x"91",x"cd"),
   781 => (x"a3",x"c1",x"81",x"f2"),
   782 => (x"c3",x"51",x"12",x"4a"),
   783 => (x"51",x"12",x"4a",x"a3"),
   784 => (x"12",x"4a",x"a3",x"c5"),
   785 => (x"4a",x"a3",x"c7",x"51"),
   786 => (x"a3",x"c9",x"51",x"12"),
   787 => (x"ce",x"51",x"12",x"4a"),
   788 => (x"51",x"12",x"4a",x"a3"),
   789 => (x"12",x"4a",x"a3",x"d0"),
   790 => (x"4a",x"a3",x"d2",x"51"),
   791 => (x"a3",x"d4",x"51",x"12"),
   792 => (x"d6",x"51",x"12",x"4a"),
   793 => (x"51",x"12",x"4a",x"a3"),
   794 => (x"12",x"4a",x"a3",x"d8"),
   795 => (x"4a",x"a3",x"dc",x"51"),
   796 => (x"a3",x"de",x"51",x"12"),
   797 => (x"c1",x"51",x"12",x"4a"),
   798 => (x"87",x"fa",x"c0",x"7e"),
   799 => (x"99",x"c8",x"49",x"74"),
   800 => (x"87",x"eb",x"c0",x"05"),
   801 => (x"99",x"d0",x"49",x"74"),
   802 => (x"dc",x"87",x"d1",x"05"),
   803 => (x"cb",x"c0",x"02",x"66"),
   804 => (x"dc",x"49",x"73",x"87"),
   805 => (x"98",x"70",x"0f",x"66"),
   806 => (x"87",x"d3",x"c0",x"02"),
   807 => (x"c6",x"c0",x"05",x"6e"),
   808 => (x"f2",x"ee",x"c2",x"87"),
   809 => (x"c0",x"50",x"c0",x"48"),
   810 => (x"48",x"bf",x"d5",x"f5"),
   811 => (x"c2",x"87",x"e1",x"c2"),
   812 => (x"c0",x"48",x"ff",x"ee"),
   813 => (x"ee",x"c2",x"7e",x"50"),
   814 => (x"c2",x"49",x"bf",x"ee"),
   815 => (x"4a",x"bf",x"de",x"e6"),
   816 => (x"fb",x"04",x"aa",x"71"),
   817 => (x"f3",x"c2",x"87",x"f6"),
   818 => (x"c0",x"05",x"bf",x"cf"),
   819 => (x"ee",x"c2",x"87",x"c8"),
   820 => (x"c1",x"02",x"bf",x"ea"),
   821 => (x"e6",x"c2",x"87",x"f8"),
   822 => (x"e9",x"49",x"bf",x"da"),
   823 => (x"49",x"70",x"87",x"c2"),
   824 => (x"59",x"de",x"e6",x"c2"),
   825 => (x"c2",x"48",x"a6",x"c4"),
   826 => (x"78",x"bf",x"da",x"e6"),
   827 => (x"bf",x"ea",x"ee",x"c2"),
   828 => (x"87",x"d8",x"c0",x"02"),
   829 => (x"cf",x"49",x"66",x"c4"),
   830 => (x"f8",x"ff",x"ff",x"ff"),
   831 => (x"c0",x"02",x"a9",x"99"),
   832 => (x"4c",x"c0",x"87",x"c5"),
   833 => (x"c1",x"87",x"e1",x"c0"),
   834 => (x"87",x"dc",x"c0",x"4c"),
   835 => (x"cf",x"49",x"66",x"c4"),
   836 => (x"a9",x"99",x"f8",x"ff"),
   837 => (x"87",x"c8",x"c0",x"02"),
   838 => (x"c0",x"48",x"a6",x"c8"),
   839 => (x"87",x"c5",x"c0",x"78"),
   840 => (x"c1",x"48",x"a6",x"c8"),
   841 => (x"4c",x"66",x"c8",x"78"),
   842 => (x"c0",x"05",x"9c",x"74"),
   843 => (x"66",x"c4",x"87",x"e0"),
   844 => (x"c2",x"89",x"c2",x"49"),
   845 => (x"4a",x"bf",x"e2",x"ee"),
   846 => (x"fb",x"f2",x"c2",x"91"),
   847 => (x"e6",x"c2",x"4a",x"bf"),
   848 => (x"a1",x"72",x"48",x"d6"),
   849 => (x"de",x"e6",x"c2",x"78"),
   850 => (x"f9",x"78",x"c0",x"48"),
   851 => (x"48",x"c0",x"87",x"de"),
   852 => (x"c3",x"e7",x"8e",x"f4"),
   853 => (x"00",x"00",x"00",x"87"),
   854 => (x"ff",x"ff",x"ff",x"00"),
   855 => (x"00",x"0d",x"65",x"ff"),
   856 => (x"00",x"0d",x"6e",x"00"),
   857 => (x"54",x"41",x"46",x"00"),
   858 => (x"20",x"20",x"32",x"33"),
   859 => (x"41",x"46",x"00",x"20"),
   860 => (x"20",x"36",x"31",x"54"),
   861 => (x"1e",x"00",x"20",x"20"),
   862 => (x"bf",x"d4",x"f3",x"c2"),
   863 => (x"05",x"a8",x"dd",x"48"),
   864 => (x"c3",x"c1",x"87",x"c9"),
   865 => (x"49",x"70",x"87",x"c8"),
   866 => (x"ff",x"87",x"c8",x"4a"),
   867 => (x"ff",x"c3",x"48",x"d4"),
   868 => (x"72",x"4a",x"68",x"78"),
   869 => (x"1e",x"4f",x"26",x"48"),
   870 => (x"bf",x"d4",x"f3",x"c2"),
   871 => (x"05",x"a8",x"dd",x"48"),
   872 => (x"c2",x"c1",x"87",x"c6"),
   873 => (x"87",x"d9",x"87",x"d4"),
   874 => (x"c3",x"48",x"d4",x"ff"),
   875 => (x"d0",x"ff",x"78",x"ff"),
   876 => (x"78",x"e1",x"c0",x"48"),
   877 => (x"d4",x"48",x"d4",x"ff"),
   878 => (x"d3",x"f3",x"c2",x"78"),
   879 => (x"bf",x"d4",x"ff",x"48"),
   880 => (x"1e",x"4f",x"26",x"50"),
   881 => (x"c0",x"48",x"d0",x"ff"),
   882 => (x"4f",x"26",x"78",x"e0"),
   883 => (x"87",x"e7",x"fe",x"1e"),
   884 => (x"02",x"99",x"49",x"70"),
   885 => (x"fb",x"c0",x"87",x"c6"),
   886 => (x"87",x"f1",x"05",x"a9"),
   887 => (x"4f",x"26",x"48",x"71"),
   888 => (x"5c",x"5b",x"5e",x"0e"),
   889 => (x"c0",x"4b",x"71",x"0e"),
   890 => (x"87",x"cb",x"fe",x"4c"),
   891 => (x"02",x"99",x"49",x"70"),
   892 => (x"c0",x"87",x"f9",x"c0"),
   893 => (x"c0",x"02",x"a9",x"ec"),
   894 => (x"fb",x"c0",x"87",x"f2"),
   895 => (x"eb",x"c0",x"02",x"a9"),
   896 => (x"b7",x"66",x"cc",x"87"),
   897 => (x"87",x"c7",x"03",x"ac"),
   898 => (x"c2",x"02",x"66",x"d0"),
   899 => (x"71",x"53",x"71",x"87"),
   900 => (x"87",x"c2",x"02",x"99"),
   901 => (x"de",x"fd",x"84",x"c1"),
   902 => (x"99",x"49",x"70",x"87"),
   903 => (x"c0",x"87",x"cd",x"02"),
   904 => (x"c7",x"02",x"a9",x"ec"),
   905 => (x"a9",x"fb",x"c0",x"87"),
   906 => (x"87",x"d5",x"ff",x"05"),
   907 => (x"c3",x"02",x"66",x"d0"),
   908 => (x"7b",x"97",x"c0",x"87"),
   909 => (x"05",x"a9",x"ec",x"c0"),
   910 => (x"4a",x"74",x"87",x"c4"),
   911 => (x"4a",x"74",x"87",x"c5"),
   912 => (x"72",x"8a",x"0a",x"c0"),
   913 => (x"26",x"87",x"c2",x"48"),
   914 => (x"26",x"4c",x"26",x"4d"),
   915 => (x"1e",x"4f",x"26",x"4b"),
   916 => (x"70",x"87",x"e4",x"fc"),
   917 => (x"b7",x"f0",x"c0",x"49"),
   918 => (x"87",x"ca",x"04",x"a9"),
   919 => (x"a9",x"b7",x"f9",x"c0"),
   920 => (x"c0",x"87",x"c3",x"01"),
   921 => (x"c1",x"c1",x"89",x"f0"),
   922 => (x"ca",x"04",x"a9",x"b7"),
   923 => (x"b7",x"da",x"c1",x"87"),
   924 => (x"87",x"c3",x"01",x"a9"),
   925 => (x"71",x"89",x"f7",x"c0"),
   926 => (x"0e",x"4f",x"26",x"48"),
   927 => (x"0e",x"5c",x"5b",x"5e"),
   928 => (x"d4",x"ff",x"4a",x"71"),
   929 => (x"c0",x"49",x"72",x"4c"),
   930 => (x"4b",x"70",x"87",x"e9"),
   931 => (x"87",x"c2",x"02",x"9b"),
   932 => (x"d0",x"ff",x"8b",x"c1"),
   933 => (x"c1",x"78",x"c5",x"48"),
   934 => (x"49",x"73",x"7c",x"d5"),
   935 => (x"e7",x"c1",x"31",x"c6"),
   936 => (x"4a",x"bf",x"97",x"d0"),
   937 => (x"70",x"b0",x"71",x"48"),
   938 => (x"48",x"d0",x"ff",x"7c"),
   939 => (x"48",x"73",x"78",x"c4"),
   940 => (x"0e",x"87",x"d6",x"fe"),
   941 => (x"5d",x"5c",x"5b",x"5e"),
   942 => (x"71",x"86",x"f4",x"0e"),
   943 => (x"48",x"a6",x"c4",x"4c"),
   944 => (x"a4",x"c8",x"78",x"c0"),
   945 => (x"bf",x"97",x"6e",x"7e"),
   946 => (x"a9",x"c1",x"c1",x"49"),
   947 => (x"c9",x"87",x"dd",x"05"),
   948 => (x"69",x"97",x"49",x"a4"),
   949 => (x"a9",x"d2",x"c1",x"49"),
   950 => (x"ca",x"87",x"d1",x"05"),
   951 => (x"69",x"97",x"49",x"a4"),
   952 => (x"a9",x"c3",x"c1",x"49"),
   953 => (x"df",x"87",x"c5",x"05"),
   954 => (x"87",x"e1",x"c2",x"48"),
   955 => (x"c0",x"87",x"e8",x"fa"),
   956 => (x"d2",x"fe",x"c0",x"4b"),
   957 => (x"c0",x"49",x"bf",x"97"),
   958 => (x"87",x"cf",x"04",x"a9"),
   959 => (x"c1",x"87",x"cd",x"fb"),
   960 => (x"d2",x"fe",x"c0",x"83"),
   961 => (x"ab",x"49",x"bf",x"97"),
   962 => (x"c0",x"87",x"f1",x"06"),
   963 => (x"bf",x"97",x"d2",x"fe"),
   964 => (x"f9",x"87",x"cf",x"02"),
   965 => (x"49",x"70",x"87",x"e1"),
   966 => (x"87",x"c6",x"02",x"99"),
   967 => (x"05",x"a9",x"ec",x"c0"),
   968 => (x"4b",x"c0",x"87",x"f1"),
   969 => (x"70",x"87",x"d0",x"f9"),
   970 => (x"87",x"cb",x"f9",x"4d"),
   971 => (x"f9",x"58",x"a6",x"cc"),
   972 => (x"4a",x"70",x"87",x"c5"),
   973 => (x"97",x"6e",x"83",x"c1"),
   974 => (x"02",x"ad",x"49",x"bf"),
   975 => (x"ff",x"c0",x"87",x"c7"),
   976 => (x"ea",x"c0",x"05",x"ad"),
   977 => (x"49",x"a4",x"c9",x"87"),
   978 => (x"c8",x"49",x"69",x"97"),
   979 => (x"c7",x"02",x"a9",x"66"),
   980 => (x"ff",x"c0",x"48",x"87"),
   981 => (x"87",x"d7",x"05",x"a8"),
   982 => (x"97",x"49",x"a4",x"ca"),
   983 => (x"02",x"aa",x"49",x"69"),
   984 => (x"ff",x"c0",x"87",x"c6"),
   985 => (x"87",x"c7",x"05",x"aa"),
   986 => (x"c1",x"48",x"a6",x"c4"),
   987 => (x"c0",x"87",x"d3",x"78"),
   988 => (x"c6",x"02",x"ad",x"ec"),
   989 => (x"ad",x"fb",x"c0",x"87"),
   990 => (x"c0",x"87",x"c7",x"05"),
   991 => (x"48",x"a6",x"c4",x"4b"),
   992 => (x"66",x"c4",x"78",x"c1"),
   993 => (x"87",x"dc",x"fe",x"02"),
   994 => (x"73",x"87",x"f8",x"f8"),
   995 => (x"fa",x"8e",x"f4",x"48"),
   996 => (x"0e",x"00",x"87",x"f5"),
   997 => (x"5d",x"5c",x"5b",x"5e"),
   998 => (x"71",x"86",x"f8",x"0e"),
   999 => (x"4b",x"d4",x"ff",x"4d"),
  1000 => (x"f3",x"c2",x"1e",x"75"),
  1001 => (x"df",x"ff",x"49",x"d8"),
  1002 => (x"86",x"c4",x"87",x"e8"),
  1003 => (x"c4",x"02",x"98",x"70"),
  1004 => (x"e7",x"c1",x"87",x"fb"),
  1005 => (x"75",x"7e",x"bf",x"d2"),
  1006 => (x"87",x"ff",x"fa",x"49"),
  1007 => (x"c0",x"05",x"a8",x"de"),
  1008 => (x"49",x"75",x"87",x"eb"),
  1009 => (x"87",x"e4",x"f7",x"c0"),
  1010 => (x"db",x"02",x"98",x"70"),
  1011 => (x"fc",x"f7",x"c2",x"87"),
  1012 => (x"e1",x"c0",x"1e",x"bf"),
  1013 => (x"cb",x"f4",x"c0",x"49"),
  1014 => (x"c1",x"86",x"c4",x"87"),
  1015 => (x"c0",x"48",x"d0",x"e7"),
  1016 => (x"c8",x"f8",x"c2",x"50"),
  1017 => (x"87",x"eb",x"fe",x"49"),
  1018 => (x"c2",x"c4",x"48",x"c1"),
  1019 => (x"48",x"d0",x"ff",x"87"),
  1020 => (x"d6",x"c1",x"78",x"c5"),
  1021 => (x"75",x"4a",x"c0",x"7b"),
  1022 => (x"7b",x"11",x"49",x"a2"),
  1023 => (x"b7",x"cb",x"82",x"c1"),
  1024 => (x"87",x"f3",x"04",x"aa"),
  1025 => (x"ff",x"c3",x"4a",x"cc"),
  1026 => (x"c0",x"82",x"c1",x"7b"),
  1027 => (x"04",x"aa",x"b7",x"e0"),
  1028 => (x"d0",x"ff",x"87",x"f4"),
  1029 => (x"c3",x"78",x"c4",x"48"),
  1030 => (x"78",x"c5",x"7b",x"ff"),
  1031 => (x"c1",x"7b",x"d3",x"c1"),
  1032 => (x"6e",x"78",x"c4",x"7b"),
  1033 => (x"a8",x"b7",x"c0",x"48"),
  1034 => (x"87",x"f0",x"c2",x"06"),
  1035 => (x"bf",x"e0",x"f3",x"c2"),
  1036 => (x"74",x"48",x"6e",x"4c"),
  1037 => (x"74",x"7e",x"70",x"88"),
  1038 => (x"fd",x"c1",x"02",x"9c"),
  1039 => (x"e2",x"e6",x"c2",x"87"),
  1040 => (x"48",x"a6",x"c4",x"4d"),
  1041 => (x"8c",x"78",x"c0",x"c8"),
  1042 => (x"03",x"ac",x"b7",x"c0"),
  1043 => (x"c0",x"c8",x"87",x"c6"),
  1044 => (x"4c",x"c0",x"78",x"a4"),
  1045 => (x"97",x"d3",x"f3",x"c2"),
  1046 => (x"99",x"d0",x"49",x"bf"),
  1047 => (x"c0",x"87",x"d1",x"02"),
  1048 => (x"d8",x"f3",x"c2",x"1e"),
  1049 => (x"87",x"dd",x"e1",x"49"),
  1050 => (x"49",x"70",x"86",x"c4"),
  1051 => (x"87",x"ee",x"c0",x"4a"),
  1052 => (x"1e",x"e2",x"e6",x"c2"),
  1053 => (x"49",x"d8",x"f3",x"c2"),
  1054 => (x"c4",x"87",x"ca",x"e1"),
  1055 => (x"4a",x"49",x"70",x"86"),
  1056 => (x"c8",x"48",x"d0",x"ff"),
  1057 => (x"d4",x"c1",x"78",x"c5"),
  1058 => (x"c4",x"7b",x"15",x"7b"),
  1059 => (x"88",x"c1",x"48",x"66"),
  1060 => (x"70",x"58",x"a6",x"c8"),
  1061 => (x"f0",x"ff",x"05",x"98"),
  1062 => (x"48",x"d0",x"ff",x"87"),
  1063 => (x"9a",x"72",x"78",x"c4"),
  1064 => (x"c0",x"87",x"c5",x"05"),
  1065 => (x"87",x"c7",x"c1",x"48"),
  1066 => (x"f3",x"c2",x"1e",x"c1"),
  1067 => (x"de",x"ff",x"49",x"d8"),
  1068 => (x"86",x"c4",x"87",x"f9"),
  1069 => (x"fe",x"05",x"9c",x"74"),
  1070 => (x"48",x"6e",x"87",x"c3"),
  1071 => (x"06",x"a8",x"b7",x"c0"),
  1072 => (x"f3",x"c2",x"87",x"d1"),
  1073 => (x"78",x"c0",x"48",x"d8"),
  1074 => (x"78",x"c0",x"80",x"d0"),
  1075 => (x"f3",x"c2",x"80",x"f4"),
  1076 => (x"6e",x"78",x"bf",x"e4"),
  1077 => (x"a8",x"b7",x"c0",x"48"),
  1078 => (x"87",x"d0",x"fd",x"01"),
  1079 => (x"c5",x"48",x"d0",x"ff"),
  1080 => (x"7b",x"d3",x"c1",x"78"),
  1081 => (x"78",x"c4",x"7b",x"c0"),
  1082 => (x"c2",x"c0",x"48",x"c1"),
  1083 => (x"f8",x"48",x"c0",x"87"),
  1084 => (x"26",x"4d",x"26",x"8e"),
  1085 => (x"26",x"4b",x"26",x"4c"),
  1086 => (x"5b",x"5e",x"0e",x"4f"),
  1087 => (x"1e",x"0e",x"5d",x"5c"),
  1088 => (x"4c",x"c0",x"4b",x"71"),
  1089 => (x"c0",x"04",x"ab",x"4d"),
  1090 => (x"fa",x"c0",x"87",x"e8"),
  1091 => (x"9d",x"75",x"1e",x"f3"),
  1092 => (x"c0",x"87",x"c4",x"02"),
  1093 => (x"c1",x"87",x"c2",x"4a"),
  1094 => (x"e9",x"49",x"72",x"4a"),
  1095 => (x"86",x"c4",x"87",x"df"),
  1096 => (x"84",x"c1",x"7e",x"70"),
  1097 => (x"87",x"c2",x"05",x"6e"),
  1098 => (x"85",x"c1",x"4c",x"73"),
  1099 => (x"ff",x"06",x"ac",x"73"),
  1100 => (x"48",x"6e",x"87",x"d8"),
  1101 => (x"87",x"f9",x"fe",x"26"),
  1102 => (x"c4",x"4a",x"71",x"1e"),
  1103 => (x"87",x"c5",x"05",x"66"),
  1104 => (x"ce",x"f9",x"49",x"72"),
  1105 => (x"0e",x"4f",x"26",x"87"),
  1106 => (x"5d",x"5c",x"5b",x"5e"),
  1107 => (x"4c",x"71",x"1e",x"0e"),
  1108 => (x"c2",x"91",x"de",x"49"),
  1109 => (x"71",x"4d",x"c0",x"f4"),
  1110 => (x"02",x"6d",x"97",x"85"),
  1111 => (x"c2",x"87",x"dc",x"c1"),
  1112 => (x"4a",x"bf",x"ec",x"f3"),
  1113 => (x"49",x"72",x"82",x"74"),
  1114 => (x"70",x"87",x"ce",x"fe"),
  1115 => (x"c0",x"02",x"6e",x"7e"),
  1116 => (x"f3",x"c2",x"87",x"f2"),
  1117 => (x"4a",x"6e",x"4b",x"f4"),
  1118 => (x"fc",x"fe",x"49",x"cb"),
  1119 => (x"4b",x"74",x"87",x"ea"),
  1120 => (x"e7",x"c1",x"93",x"cb"),
  1121 => (x"83",x"c4",x"83",x"e4"),
  1122 => (x"7b",x"ff",x"c6",x"c1"),
  1123 => (x"cc",x"c1",x"49",x"74"),
  1124 => (x"7b",x"75",x"87",x"c7"),
  1125 => (x"97",x"d1",x"e7",x"c1"),
  1126 => (x"c2",x"1e",x"49",x"bf"),
  1127 => (x"fe",x"49",x"f4",x"f3"),
  1128 => (x"86",x"c4",x"87",x"d6"),
  1129 => (x"cb",x"c1",x"49",x"74"),
  1130 => (x"49",x"c0",x"87",x"ef"),
  1131 => (x"87",x"ce",x"cd",x"c1"),
  1132 => (x"48",x"d4",x"f3",x"c2"),
  1133 => (x"49",x"c1",x"78",x"c0"),
  1134 => (x"26",x"87",x"d4",x"dd"),
  1135 => (x"4c",x"87",x"f2",x"fc"),
  1136 => (x"69",x"64",x"61",x"6f"),
  1137 => (x"2e",x"2e",x"67",x"6e"),
  1138 => (x"5e",x"0e",x"00",x"2e"),
  1139 => (x"71",x"0e",x"5c",x"5b"),
  1140 => (x"f3",x"c2",x"4a",x"4b"),
  1141 => (x"72",x"82",x"bf",x"ec"),
  1142 => (x"87",x"dd",x"fc",x"49"),
  1143 => (x"02",x"9c",x"4c",x"70"),
  1144 => (x"e5",x"49",x"87",x"c4"),
  1145 => (x"f3",x"c2",x"87",x"df"),
  1146 => (x"78",x"c0",x"48",x"ec"),
  1147 => (x"de",x"dc",x"49",x"c1"),
  1148 => (x"87",x"ff",x"fb",x"87"),
  1149 => (x"5c",x"5b",x"5e",x"0e"),
  1150 => (x"86",x"f4",x"0e",x"5d"),
  1151 => (x"4d",x"e2",x"e6",x"c2"),
  1152 => (x"a6",x"c4",x"4c",x"c0"),
  1153 => (x"c2",x"78",x"c0",x"48"),
  1154 => (x"49",x"bf",x"ec",x"f3"),
  1155 => (x"c1",x"06",x"a9",x"c0"),
  1156 => (x"e6",x"c2",x"87",x"c1"),
  1157 => (x"02",x"98",x"48",x"e2"),
  1158 => (x"c0",x"87",x"f8",x"c0"),
  1159 => (x"c8",x"1e",x"f3",x"fa"),
  1160 => (x"87",x"c7",x"02",x"66"),
  1161 => (x"c0",x"48",x"a6",x"c4"),
  1162 => (x"c4",x"87",x"c5",x"78"),
  1163 => (x"78",x"c1",x"48",x"a6"),
  1164 => (x"e5",x"49",x"66",x"c4"),
  1165 => (x"86",x"c4",x"87",x"c7"),
  1166 => (x"84",x"c1",x"4d",x"70"),
  1167 => (x"c1",x"48",x"66",x"c4"),
  1168 => (x"58",x"a6",x"c8",x"80"),
  1169 => (x"bf",x"ec",x"f3",x"c2"),
  1170 => (x"c6",x"03",x"ac",x"49"),
  1171 => (x"05",x"9d",x"75",x"87"),
  1172 => (x"c0",x"87",x"c8",x"ff"),
  1173 => (x"02",x"9d",x"75",x"4c"),
  1174 => (x"c0",x"87",x"e0",x"c3"),
  1175 => (x"c8",x"1e",x"f3",x"fa"),
  1176 => (x"87",x"c7",x"02",x"66"),
  1177 => (x"c0",x"48",x"a6",x"cc"),
  1178 => (x"cc",x"87",x"c5",x"78"),
  1179 => (x"78",x"c1",x"48",x"a6"),
  1180 => (x"e4",x"49",x"66",x"cc"),
  1181 => (x"86",x"c4",x"87",x"c7"),
  1182 => (x"02",x"6e",x"7e",x"70"),
  1183 => (x"6e",x"87",x"e9",x"c2"),
  1184 => (x"97",x"81",x"cb",x"49"),
  1185 => (x"99",x"d0",x"49",x"69"),
  1186 => (x"87",x"d6",x"c1",x"02"),
  1187 => (x"4a",x"ca",x"c7",x"c1"),
  1188 => (x"91",x"cb",x"49",x"74"),
  1189 => (x"81",x"e4",x"e7",x"c1"),
  1190 => (x"81",x"c8",x"79",x"72"),
  1191 => (x"74",x"51",x"ff",x"c3"),
  1192 => (x"c2",x"91",x"de",x"49"),
  1193 => (x"71",x"4d",x"c0",x"f4"),
  1194 => (x"97",x"c1",x"c2",x"85"),
  1195 => (x"49",x"a5",x"c1",x"7d"),
  1196 => (x"c2",x"51",x"e0",x"c0"),
  1197 => (x"bf",x"97",x"f2",x"ee"),
  1198 => (x"c1",x"87",x"d2",x"02"),
  1199 => (x"4b",x"a5",x"c2",x"84"),
  1200 => (x"4a",x"f2",x"ee",x"c2"),
  1201 => (x"f7",x"fe",x"49",x"db"),
  1202 => (x"db",x"c1",x"87",x"de"),
  1203 => (x"49",x"a5",x"cd",x"87"),
  1204 => (x"84",x"c1",x"51",x"c0"),
  1205 => (x"6e",x"4b",x"a5",x"c2"),
  1206 => (x"fe",x"49",x"cb",x"4a"),
  1207 => (x"c1",x"87",x"c9",x"f7"),
  1208 => (x"c5",x"c1",x"87",x"c6"),
  1209 => (x"49",x"74",x"4a",x"c7"),
  1210 => (x"e7",x"c1",x"91",x"cb"),
  1211 => (x"79",x"72",x"81",x"e4"),
  1212 => (x"97",x"f2",x"ee",x"c2"),
  1213 => (x"87",x"d8",x"02",x"bf"),
  1214 => (x"91",x"de",x"49",x"74"),
  1215 => (x"f4",x"c2",x"84",x"c1"),
  1216 => (x"83",x"71",x"4b",x"c0"),
  1217 => (x"4a",x"f2",x"ee",x"c2"),
  1218 => (x"f6",x"fe",x"49",x"dd"),
  1219 => (x"87",x"d8",x"87",x"da"),
  1220 => (x"93",x"de",x"4b",x"74"),
  1221 => (x"83",x"c0",x"f4",x"c2"),
  1222 => (x"c0",x"49",x"a3",x"cb"),
  1223 => (x"73",x"84",x"c1",x"51"),
  1224 => (x"49",x"cb",x"4a",x"6e"),
  1225 => (x"87",x"c0",x"f6",x"fe"),
  1226 => (x"c1",x"48",x"66",x"c4"),
  1227 => (x"58",x"a6",x"c8",x"80"),
  1228 => (x"c0",x"03",x"ac",x"c7"),
  1229 => (x"05",x"6e",x"87",x"c5"),
  1230 => (x"74",x"87",x"e0",x"fc"),
  1231 => (x"f6",x"8e",x"f4",x"48"),
  1232 => (x"73",x"1e",x"87",x"ef"),
  1233 => (x"49",x"4b",x"71",x"1e"),
  1234 => (x"e7",x"c1",x"91",x"cb"),
  1235 => (x"a1",x"c8",x"81",x"e4"),
  1236 => (x"d0",x"e7",x"c1",x"4a"),
  1237 => (x"c9",x"50",x"12",x"48"),
  1238 => (x"fe",x"c0",x"4a",x"a1"),
  1239 => (x"50",x"12",x"48",x"d2"),
  1240 => (x"e7",x"c1",x"81",x"ca"),
  1241 => (x"50",x"11",x"48",x"d1"),
  1242 => (x"97",x"d1",x"e7",x"c1"),
  1243 => (x"c0",x"1e",x"49",x"bf"),
  1244 => (x"87",x"c4",x"f7",x"49"),
  1245 => (x"48",x"d4",x"f3",x"c2"),
  1246 => (x"49",x"c1",x"78",x"de"),
  1247 => (x"26",x"87",x"d0",x"d6"),
  1248 => (x"1e",x"87",x"f2",x"f5"),
  1249 => (x"cb",x"49",x"4a",x"71"),
  1250 => (x"e4",x"e7",x"c1",x"91"),
  1251 => (x"11",x"81",x"c8",x"81"),
  1252 => (x"d8",x"f3",x"c2",x"48"),
  1253 => (x"ec",x"f3",x"c2",x"58"),
  1254 => (x"c1",x"78",x"c0",x"48"),
  1255 => (x"87",x"ef",x"d5",x"49"),
  1256 => (x"c0",x"1e",x"4f",x"26"),
  1257 => (x"d5",x"c5",x"c1",x"49"),
  1258 => (x"1e",x"4f",x"26",x"87"),
  1259 => (x"d2",x"02",x"99",x"71"),
  1260 => (x"f9",x"e8",x"c1",x"87"),
  1261 => (x"f7",x"50",x"c0",x"48"),
  1262 => (x"c3",x"ce",x"c1",x"80"),
  1263 => (x"dd",x"e7",x"c1",x"40"),
  1264 => (x"c1",x"87",x"ce",x"78"),
  1265 => (x"c1",x"48",x"f5",x"e8"),
  1266 => (x"fc",x"78",x"d6",x"e7"),
  1267 => (x"e2",x"ce",x"c1",x"80"),
  1268 => (x"0e",x"4f",x"26",x"78"),
  1269 => (x"0e",x"5c",x"5b",x"5e"),
  1270 => (x"cb",x"4a",x"4c",x"71"),
  1271 => (x"e4",x"e7",x"c1",x"92"),
  1272 => (x"49",x"a2",x"c8",x"82"),
  1273 => (x"97",x"4b",x"a2",x"c9"),
  1274 => (x"97",x"1e",x"4b",x"6b"),
  1275 => (x"ca",x"1e",x"49",x"69"),
  1276 => (x"c0",x"49",x"12",x"82"),
  1277 => (x"c0",x"87",x"f5",x"e5"),
  1278 => (x"87",x"d3",x"d4",x"49"),
  1279 => (x"c2",x"c1",x"49",x"74"),
  1280 => (x"8e",x"f8",x"87",x"d7"),
  1281 => (x"1e",x"87",x"ec",x"f3"),
  1282 => (x"4b",x"71",x"1e",x"73"),
  1283 => (x"87",x"c3",x"ff",x"49"),
  1284 => (x"fe",x"fe",x"49",x"73"),
  1285 => (x"87",x"dd",x"f3",x"87"),
  1286 => (x"71",x"1e",x"73",x"1e"),
  1287 => (x"4a",x"a3",x"c6",x"4b"),
  1288 => (x"c1",x"87",x"db",x"02"),
  1289 => (x"87",x"d6",x"02",x"8a"),
  1290 => (x"da",x"c1",x"02",x"8a"),
  1291 => (x"c0",x"02",x"8a",x"87"),
  1292 => (x"02",x"8a",x"87",x"fc"),
  1293 => (x"8a",x"87",x"e1",x"c0"),
  1294 => (x"c1",x"87",x"cb",x"02"),
  1295 => (x"49",x"c7",x"87",x"db"),
  1296 => (x"c1",x"87",x"c0",x"fd"),
  1297 => (x"f3",x"c2",x"87",x"de"),
  1298 => (x"c1",x"02",x"bf",x"ec"),
  1299 => (x"c1",x"48",x"87",x"cb"),
  1300 => (x"f0",x"f3",x"c2",x"88"),
  1301 => (x"87",x"c1",x"c1",x"58"),
  1302 => (x"bf",x"f0",x"f3",x"c2"),
  1303 => (x"87",x"f9",x"c0",x"02"),
  1304 => (x"bf",x"ec",x"f3",x"c2"),
  1305 => (x"c2",x"80",x"c1",x"48"),
  1306 => (x"c0",x"58",x"f0",x"f3"),
  1307 => (x"f3",x"c2",x"87",x"eb"),
  1308 => (x"c6",x"49",x"bf",x"ec"),
  1309 => (x"f0",x"f3",x"c2",x"89"),
  1310 => (x"a9",x"b7",x"c0",x"59"),
  1311 => (x"c2",x"87",x"da",x"03"),
  1312 => (x"c0",x"48",x"ec",x"f3"),
  1313 => (x"c2",x"87",x"d2",x"78"),
  1314 => (x"02",x"bf",x"f0",x"f3"),
  1315 => (x"f3",x"c2",x"87",x"cb"),
  1316 => (x"c6",x"48",x"bf",x"ec"),
  1317 => (x"f0",x"f3",x"c2",x"80"),
  1318 => (x"d1",x"49",x"c0",x"58"),
  1319 => (x"49",x"73",x"87",x"f1"),
  1320 => (x"87",x"f5",x"ff",x"c0"),
  1321 => (x"1e",x"87",x"ce",x"f1"),
  1322 => (x"4b",x"71",x"1e",x"73"),
  1323 => (x"48",x"d4",x"f3",x"c2"),
  1324 => (x"49",x"c0",x"78",x"dd"),
  1325 => (x"73",x"87",x"d8",x"d1"),
  1326 => (x"dc",x"ff",x"c0",x"49"),
  1327 => (x"87",x"f5",x"f0",x"87"),
  1328 => (x"5c",x"5b",x"5e",x"0e"),
  1329 => (x"cc",x"4c",x"71",x"0e"),
  1330 => (x"4b",x"74",x"1e",x"66"),
  1331 => (x"e7",x"c1",x"93",x"cb"),
  1332 => (x"a3",x"c4",x"83",x"e4"),
  1333 => (x"fe",x"49",x"6a",x"4a"),
  1334 => (x"c1",x"87",x"dd",x"ef"),
  1335 => (x"c8",x"7b",x"c2",x"cd"),
  1336 => (x"66",x"d4",x"49",x"a3"),
  1337 => (x"49",x"a3",x"c9",x"51"),
  1338 => (x"ca",x"51",x"66",x"d8"),
  1339 => (x"66",x"dc",x"49",x"a3"),
  1340 => (x"fe",x"ef",x"26",x"51"),
  1341 => (x"5b",x"5e",x"0e",x"87"),
  1342 => (x"ff",x"0e",x"5d",x"5c"),
  1343 => (x"a6",x"dc",x"86",x"cc"),
  1344 => (x"48",x"a6",x"c8",x"59"),
  1345 => (x"80",x"c4",x"78",x"c0"),
  1346 => (x"78",x"66",x"c8",x"c1"),
  1347 => (x"78",x"c1",x"80",x"c4"),
  1348 => (x"78",x"c1",x"80",x"c4"),
  1349 => (x"48",x"f0",x"f3",x"c2"),
  1350 => (x"f3",x"c2",x"78",x"c1"),
  1351 => (x"de",x"48",x"bf",x"d4"),
  1352 => (x"87",x"cb",x"05",x"a8"),
  1353 => (x"70",x"87",x"cd",x"f3"),
  1354 => (x"59",x"a6",x"cc",x"49"),
  1355 => (x"e1",x"87",x"db",x"ce"),
  1356 => (x"d7",x"e2",x"87",x"e5"),
  1357 => (x"87",x"ff",x"e0",x"87"),
  1358 => (x"fb",x"c0",x"4c",x"70"),
  1359 => (x"dd",x"c1",x"02",x"ac"),
  1360 => (x"05",x"66",x"d8",x"87"),
  1361 => (x"c0",x"87",x"cf",x"c1"),
  1362 => (x"1e",x"c1",x"1e",x"1e"),
  1363 => (x"1e",x"c7",x"e9",x"c1"),
  1364 => (x"eb",x"fd",x"49",x"c0"),
  1365 => (x"c1",x"86",x"d0",x"87"),
  1366 => (x"c4",x"48",x"66",x"c4"),
  1367 => (x"6e",x"7e",x"70",x"80"),
  1368 => (x"81",x"c7",x"49",x"bf"),
  1369 => (x"fb",x"c0",x"51",x"74"),
  1370 => (x"87",x"cf",x"02",x"ac"),
  1371 => (x"1e",x"d8",x"1e",x"c1"),
  1372 => (x"49",x"bf",x"66",x"c8"),
  1373 => (x"e7",x"e1",x"81",x"c8"),
  1374 => (x"c1",x"86",x"c8",x"87"),
  1375 => (x"c0",x"48",x"66",x"c8"),
  1376 => (x"87",x"c7",x"01",x"a8"),
  1377 => (x"c1",x"48",x"a6",x"c8"),
  1378 => (x"c1",x"87",x"ce",x"78"),
  1379 => (x"c1",x"48",x"66",x"c8"),
  1380 => (x"58",x"a6",x"d0",x"88"),
  1381 => (x"f3",x"e0",x"87",x"c3"),
  1382 => (x"48",x"a6",x"d0",x"87"),
  1383 => (x"9c",x"74",x"78",x"c2"),
  1384 => (x"87",x"e2",x"cc",x"02"),
  1385 => (x"c1",x"48",x"66",x"c8"),
  1386 => (x"03",x"a8",x"66",x"cc"),
  1387 => (x"c4",x"87",x"d7",x"cc"),
  1388 => (x"78",x"c0",x"48",x"a6"),
  1389 => (x"78",x"c0",x"80",x"d8"),
  1390 => (x"87",x"fb",x"de",x"ff"),
  1391 => (x"66",x"d8",x"4c",x"70"),
  1392 => (x"05",x"a8",x"dd",x"48"),
  1393 => (x"a6",x"dc",x"87",x"c6"),
  1394 => (x"78",x"66",x"d8",x"48"),
  1395 => (x"05",x"ac",x"d0",x"c1"),
  1396 => (x"ff",x"87",x"eb",x"c0"),
  1397 => (x"ff",x"87",x"e0",x"de"),
  1398 => (x"70",x"87",x"dc",x"de"),
  1399 => (x"ac",x"ec",x"c0",x"4c"),
  1400 => (x"ff",x"87",x"c6",x"05"),
  1401 => (x"70",x"87",x"e5",x"df"),
  1402 => (x"ac",x"d0",x"c1",x"4c"),
  1403 => (x"d4",x"87",x"c8",x"05"),
  1404 => (x"80",x"c1",x"48",x"66"),
  1405 => (x"c1",x"58",x"a6",x"d8"),
  1406 => (x"ff",x"02",x"ac",x"d0"),
  1407 => (x"e0",x"c0",x"87",x"d5"),
  1408 => (x"66",x"d8",x"48",x"a6"),
  1409 => (x"48",x"66",x"dc",x"78"),
  1410 => (x"a8",x"66",x"e0",x"c0"),
  1411 => (x"87",x"c8",x"ca",x"05"),
  1412 => (x"48",x"a6",x"e4",x"c0"),
  1413 => (x"80",x"c4",x"78",x"c0"),
  1414 => (x"4d",x"74",x"78",x"c0"),
  1415 => (x"02",x"8d",x"fb",x"c0"),
  1416 => (x"c9",x"87",x"ce",x"c9"),
  1417 => (x"87",x"db",x"02",x"8d"),
  1418 => (x"c1",x"02",x"8d",x"c2"),
  1419 => (x"8d",x"c9",x"87",x"f7"),
  1420 => (x"87",x"d1",x"c4",x"02"),
  1421 => (x"c1",x"02",x"8d",x"c4"),
  1422 => (x"8d",x"c1",x"87",x"c2"),
  1423 => (x"87",x"c5",x"c4",x"02"),
  1424 => (x"c8",x"87",x"e8",x"c8"),
  1425 => (x"91",x"cb",x"49",x"66"),
  1426 => (x"81",x"66",x"c4",x"c1"),
  1427 => (x"6a",x"4a",x"a1",x"c4"),
  1428 => (x"c1",x"1e",x"71",x"7e"),
  1429 => (x"c4",x"48",x"c2",x"e4"),
  1430 => (x"a1",x"cc",x"49",x"66"),
  1431 => (x"71",x"41",x"20",x"4a"),
  1432 => (x"f8",x"ff",x"05",x"aa"),
  1433 => (x"26",x"51",x"10",x"87"),
  1434 => (x"e7",x"d2",x"c1",x"49"),
  1435 => (x"db",x"dd",x"ff",x"79"),
  1436 => (x"c0",x"4c",x"70",x"87"),
  1437 => (x"c1",x"48",x"a6",x"e8"),
  1438 => (x"87",x"f5",x"c7",x"78"),
  1439 => (x"c0",x"48",x"a6",x"c4"),
  1440 => (x"db",x"ff",x"78",x"f0"),
  1441 => (x"4c",x"70",x"87",x"f1"),
  1442 => (x"02",x"ac",x"ec",x"c0"),
  1443 => (x"c8",x"87",x"c3",x"c0"),
  1444 => (x"ec",x"c0",x"5c",x"a6"),
  1445 => (x"87",x"cd",x"02",x"ac"),
  1446 => (x"87",x"db",x"db",x"ff"),
  1447 => (x"ec",x"c0",x"4c",x"70"),
  1448 => (x"f3",x"ff",x"05",x"ac"),
  1449 => (x"ac",x"ec",x"c0",x"87"),
  1450 => (x"87",x"c4",x"c0",x"02"),
  1451 => (x"87",x"c7",x"db",x"ff"),
  1452 => (x"d8",x"1e",x"66",x"c4"),
  1453 => (x"d8",x"1e",x"49",x"66"),
  1454 => (x"c1",x"1e",x"49",x"66"),
  1455 => (x"d8",x"1e",x"c7",x"e9"),
  1456 => (x"fb",x"f7",x"49",x"66"),
  1457 => (x"ca",x"1e",x"c0",x"87"),
  1458 => (x"66",x"e0",x"c0",x"1e"),
  1459 => (x"c1",x"91",x"cb",x"49"),
  1460 => (x"d8",x"81",x"66",x"dc"),
  1461 => (x"a1",x"c4",x"48",x"a6"),
  1462 => (x"bf",x"66",x"d8",x"78"),
  1463 => (x"ff",x"db",x"ff",x"49"),
  1464 => (x"c0",x"86",x"d8",x"87"),
  1465 => (x"c1",x"06",x"a8",x"b7"),
  1466 => (x"1e",x"c1",x"87",x"cb"),
  1467 => (x"66",x"c8",x"1e",x"de"),
  1468 => (x"db",x"ff",x"49",x"bf"),
  1469 => (x"86",x"c8",x"87",x"ea"),
  1470 => (x"c0",x"48",x"49",x"70"),
  1471 => (x"ec",x"c0",x"88",x"08"),
  1472 => (x"b7",x"c0",x"58",x"a6"),
  1473 => (x"ec",x"c0",x"06",x"a8"),
  1474 => (x"66",x"e8",x"c0",x"87"),
  1475 => (x"a8",x"b7",x"dd",x"48"),
  1476 => (x"87",x"e1",x"c0",x"03"),
  1477 => (x"c0",x"49",x"bf",x"6e"),
  1478 => (x"c0",x"81",x"66",x"e8"),
  1479 => (x"e8",x"c0",x"51",x"e0"),
  1480 => (x"81",x"c1",x"49",x"66"),
  1481 => (x"c2",x"81",x"bf",x"6e"),
  1482 => (x"e8",x"c0",x"51",x"c1"),
  1483 => (x"81",x"c2",x"49",x"66"),
  1484 => (x"c0",x"81",x"bf",x"6e"),
  1485 => (x"48",x"66",x"d0",x"51"),
  1486 => (x"a6",x"d4",x"80",x"c1"),
  1487 => (x"80",x"d8",x"48",x"58"),
  1488 => (x"ec",x"c4",x"78",x"c1"),
  1489 => (x"c6",x"dc",x"ff",x"87"),
  1490 => (x"a6",x"ec",x"c0",x"87"),
  1491 => (x"fe",x"db",x"ff",x"58"),
  1492 => (x"a6",x"f0",x"c0",x"87"),
  1493 => (x"a8",x"ec",x"c0",x"58"),
  1494 => (x"87",x"c9",x"c0",x"05"),
  1495 => (x"e8",x"c0",x"48",x"a6"),
  1496 => (x"c4",x"c0",x"78",x"66"),
  1497 => (x"ce",x"d8",x"ff",x"87"),
  1498 => (x"49",x"66",x"c8",x"87"),
  1499 => (x"c4",x"c1",x"91",x"cb"),
  1500 => (x"80",x"71",x"48",x"66"),
  1501 => (x"c4",x"58",x"a6",x"c8"),
  1502 => (x"82",x"c8",x"4a",x"66"),
  1503 => (x"ca",x"49",x"66",x"c4"),
  1504 => (x"66",x"e8",x"c0",x"81"),
  1505 => (x"66",x"ec",x"c0",x"51"),
  1506 => (x"c0",x"81",x"c1",x"49"),
  1507 => (x"c1",x"89",x"66",x"e8"),
  1508 => (x"70",x"30",x"71",x"48"),
  1509 => (x"71",x"89",x"c1",x"49"),
  1510 => (x"f7",x"c2",x"7a",x"97"),
  1511 => (x"c0",x"49",x"bf",x"dc"),
  1512 => (x"97",x"29",x"66",x"e8"),
  1513 => (x"71",x"48",x"4a",x"6a"),
  1514 => (x"a6",x"f4",x"c0",x"98"),
  1515 => (x"49",x"66",x"c4",x"58"),
  1516 => (x"7e",x"69",x"81",x"c4"),
  1517 => (x"48",x"66",x"e0",x"c0"),
  1518 => (x"02",x"a8",x"66",x"dc"),
  1519 => (x"dc",x"87",x"c8",x"c0"),
  1520 => (x"78",x"c0",x"48",x"a6"),
  1521 => (x"dc",x"87",x"c5",x"c0"),
  1522 => (x"78",x"c1",x"48",x"a6"),
  1523 => (x"c0",x"1e",x"66",x"dc"),
  1524 => (x"66",x"c8",x"1e",x"e0"),
  1525 => (x"c7",x"d8",x"ff",x"49"),
  1526 => (x"70",x"86",x"c8",x"87"),
  1527 => (x"ac",x"b7",x"c0",x"4c"),
  1528 => (x"87",x"d6",x"c1",x"06"),
  1529 => (x"80",x"74",x"48",x"6e"),
  1530 => (x"e0",x"c0",x"7e",x"70"),
  1531 => (x"6e",x"89",x"74",x"49"),
  1532 => (x"ff",x"e3",x"c1",x"4b"),
  1533 => (x"e2",x"fe",x"71",x"4a"),
  1534 => (x"48",x"6e",x"87",x"ee"),
  1535 => (x"7e",x"70",x"80",x"c2"),
  1536 => (x"48",x"66",x"e4",x"c0"),
  1537 => (x"e8",x"c0",x"80",x"c1"),
  1538 => (x"f0",x"c0",x"58",x"a6"),
  1539 => (x"81",x"c1",x"49",x"66"),
  1540 => (x"c0",x"02",x"a9",x"70"),
  1541 => (x"4d",x"c0",x"87",x"c5"),
  1542 => (x"c1",x"87",x"c2",x"c0"),
  1543 => (x"c2",x"1e",x"75",x"4d"),
  1544 => (x"e0",x"c0",x"49",x"a4"),
  1545 => (x"70",x"88",x"71",x"48"),
  1546 => (x"66",x"c8",x"1e",x"49"),
  1547 => (x"ef",x"d6",x"ff",x"49"),
  1548 => (x"c0",x"86",x"c8",x"87"),
  1549 => (x"ff",x"01",x"a8",x"b7"),
  1550 => (x"e4",x"c0",x"87",x"c6"),
  1551 => (x"d3",x"c0",x"02",x"66"),
  1552 => (x"49",x"66",x"c4",x"87"),
  1553 => (x"e4",x"c0",x"81",x"c9"),
  1554 => (x"66",x"c4",x"51",x"66"),
  1555 => (x"d3",x"cf",x"c1",x"48"),
  1556 => (x"87",x"ce",x"c0",x"78"),
  1557 => (x"c9",x"49",x"66",x"c4"),
  1558 => (x"c4",x"51",x"c2",x"81"),
  1559 => (x"d0",x"c1",x"48",x"66"),
  1560 => (x"e8",x"c0",x"78",x"c7"),
  1561 => (x"78",x"c1",x"48",x"a6"),
  1562 => (x"ff",x"87",x"c6",x"c0"),
  1563 => (x"70",x"87",x"dd",x"d5"),
  1564 => (x"66",x"e8",x"c0",x"4c"),
  1565 => (x"87",x"f5",x"c0",x"02"),
  1566 => (x"cc",x"48",x"66",x"c8"),
  1567 => (x"c0",x"04",x"a8",x"66"),
  1568 => (x"66",x"c8",x"87",x"cb"),
  1569 => (x"cc",x"80",x"c1",x"48"),
  1570 => (x"e0",x"c0",x"58",x"a6"),
  1571 => (x"48",x"66",x"cc",x"87"),
  1572 => (x"a6",x"d0",x"88",x"c1"),
  1573 => (x"87",x"d5",x"c0",x"58"),
  1574 => (x"05",x"ac",x"c6",x"c1"),
  1575 => (x"d0",x"87",x"c8",x"c0"),
  1576 => (x"80",x"c1",x"48",x"66"),
  1577 => (x"ff",x"58",x"a6",x"d4"),
  1578 => (x"70",x"87",x"e1",x"d4"),
  1579 => (x"48",x"66",x"d4",x"4c"),
  1580 => (x"a6",x"d8",x"80",x"c1"),
  1581 => (x"02",x"9c",x"74",x"58"),
  1582 => (x"c8",x"87",x"cb",x"c0"),
  1583 => (x"cc",x"c1",x"48",x"66"),
  1584 => (x"f3",x"04",x"a8",x"66"),
  1585 => (x"d3",x"ff",x"87",x"e9"),
  1586 => (x"66",x"c8",x"87",x"f9"),
  1587 => (x"03",x"a8",x"c7",x"48"),
  1588 => (x"c2",x"87",x"e5",x"c0"),
  1589 => (x"c0",x"48",x"f0",x"f3"),
  1590 => (x"49",x"66",x"c8",x"78"),
  1591 => (x"c4",x"c1",x"91",x"cb"),
  1592 => (x"a1",x"c4",x"81",x"66"),
  1593 => (x"c0",x"4a",x"6a",x"4a"),
  1594 => (x"66",x"c8",x"79",x"52"),
  1595 => (x"cc",x"80",x"c1",x"48"),
  1596 => (x"a8",x"c7",x"58",x"a6"),
  1597 => (x"87",x"db",x"ff",x"04"),
  1598 => (x"ff",x"8e",x"cc",x"ff"),
  1599 => (x"3a",x"87",x"f2",x"df"),
  1600 => (x"49",x"44",x"00",x"20"),
  1601 => (x"77",x"53",x"20",x"50"),
  1602 => (x"68",x"63",x"74",x"69"),
  1603 => (x"1e",x"00",x"73",x"65"),
  1604 => (x"4b",x"71",x"1e",x"73"),
  1605 => (x"87",x"c6",x"02",x"9b"),
  1606 => (x"48",x"ec",x"f3",x"c2"),
  1607 => (x"1e",x"c7",x"78",x"c0"),
  1608 => (x"bf",x"ec",x"f3",x"c2"),
  1609 => (x"e7",x"c1",x"1e",x"49"),
  1610 => (x"f3",x"c2",x"1e",x"e4"),
  1611 => (x"ef",x"49",x"bf",x"d4"),
  1612 => (x"86",x"cc",x"87",x"c3"),
  1613 => (x"bf",x"d4",x"f3",x"c2"),
  1614 => (x"87",x"ef",x"e9",x"49"),
  1615 => (x"c8",x"02",x"9b",x"73"),
  1616 => (x"e4",x"e7",x"c1",x"87"),
  1617 => (x"e2",x"ee",x"c0",x"49"),
  1618 => (x"e8",x"de",x"ff",x"87"),
  1619 => (x"d5",x"c7",x"1e",x"87"),
  1620 => (x"fe",x"49",x"c1",x"87"),
  1621 => (x"e5",x"fe",x"87",x"f9"),
  1622 => (x"98",x"70",x"87",x"e9"),
  1623 => (x"fe",x"87",x"cd",x"02"),
  1624 => (x"70",x"87",x"c2",x"ed"),
  1625 => (x"87",x"c4",x"02",x"98"),
  1626 => (x"87",x"c2",x"4a",x"c1"),
  1627 => (x"9a",x"72",x"4a",x"c0"),
  1628 => (x"c0",x"87",x"ce",x"05"),
  1629 => (x"e2",x"e6",x"c1",x"1e"),
  1630 => (x"cc",x"fa",x"c0",x"49"),
  1631 => (x"fe",x"86",x"c4",x"87"),
  1632 => (x"ef",x"fc",x"c0",x"87"),
  1633 => (x"c1",x"1e",x"c0",x"87"),
  1634 => (x"c0",x"49",x"ed",x"e6"),
  1635 => (x"c0",x"87",x"fa",x"f9"),
  1636 => (x"f5",x"fe",x"c0",x"1e"),
  1637 => (x"c0",x"49",x"70",x"87"),
  1638 => (x"c3",x"87",x"ee",x"f9"),
  1639 => (x"8e",x"f8",x"87",x"c7"),
  1640 => (x"44",x"53",x"4f",x"26"),
  1641 => (x"69",x"61",x"66",x"20"),
  1642 => (x"2e",x"64",x"65",x"6c"),
  1643 => (x"6f",x"6f",x"42",x"00"),
  1644 => (x"67",x"6e",x"69",x"74"),
  1645 => (x"00",x"2e",x"2e",x"2e"),
  1646 => (x"ec",x"f3",x"c2",x"1e"),
  1647 => (x"c2",x"78",x"c0",x"48"),
  1648 => (x"c0",x"48",x"d4",x"f3"),
  1649 => (x"87",x"c5",x"fe",x"78"),
  1650 => (x"87",x"dd",x"fe",x"c0"),
  1651 => (x"4f",x"26",x"48",x"c0"),
  1652 => (x"00",x"01",x"00",x"00"),
  1653 => (x"20",x"80",x"00",x"00"),
  1654 => (x"74",x"69",x"78",x"45"),
  1655 => (x"42",x"20",x"80",x"00"),
  1656 => (x"00",x"6b",x"63",x"61"),
  1657 => (x"00",x"00",x"13",x"83"),
  1658 => (x"00",x"00",x"2d",x"00"),
  1659 => (x"83",x"00",x"00",x"00"),
  1660 => (x"1e",x"00",x"00",x"13"),
  1661 => (x"00",x"00",x"00",x"2d"),
  1662 => (x"13",x"83",x"00",x"00"),
  1663 => (x"2d",x"3c",x"00",x"00"),
  1664 => (x"00",x"00",x"00",x"00"),
  1665 => (x"00",x"13",x"83",x"00"),
  1666 => (x"00",x"2d",x"5a",x"00"),
  1667 => (x"00",x"00",x"00",x"00"),
  1668 => (x"00",x"00",x"13",x"83"),
  1669 => (x"00",x"00",x"2d",x"78"),
  1670 => (x"83",x"00",x"00",x"00"),
  1671 => (x"96",x"00",x"00",x"13"),
  1672 => (x"00",x"00",x"00",x"2d"),
  1673 => (x"13",x"83",x"00",x"00"),
  1674 => (x"2d",x"b4",x"00",x"00"),
  1675 => (x"00",x"00",x"00",x"00"),
  1676 => (x"00",x"13",x"83",x"00"),
  1677 => (x"00",x"00",x"00",x"00"),
  1678 => (x"00",x"00",x"00",x"00"),
  1679 => (x"00",x"00",x"14",x"18"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"4c",x"00",x"00",x"00"),
  1682 => (x"20",x"64",x"61",x"6f"),
  1683 => (x"1e",x"00",x"2e",x"2a"),
  1684 => (x"c0",x"48",x"f0",x"fe"),
  1685 => (x"79",x"09",x"cd",x"78"),
  1686 => (x"1e",x"4f",x"26",x"09"),
  1687 => (x"bf",x"f0",x"fe",x"1e"),
  1688 => (x"26",x"26",x"48",x"7e"),
  1689 => (x"f0",x"fe",x"1e",x"4f"),
  1690 => (x"26",x"78",x"c1",x"48"),
  1691 => (x"f0",x"fe",x"1e",x"4f"),
  1692 => (x"26",x"78",x"c0",x"48"),
  1693 => (x"4a",x"71",x"1e",x"4f"),
  1694 => (x"26",x"52",x"52",x"c0"),
  1695 => (x"5b",x"5e",x"0e",x"4f"),
  1696 => (x"f4",x"0e",x"5d",x"5c"),
  1697 => (x"97",x"4d",x"71",x"86"),
  1698 => (x"a5",x"c1",x"7e",x"6d"),
  1699 => (x"48",x"6c",x"97",x"4c"),
  1700 => (x"6e",x"58",x"a6",x"c8"),
  1701 => (x"a8",x"66",x"c4",x"48"),
  1702 => (x"ff",x"87",x"c5",x"05"),
  1703 => (x"87",x"e6",x"c0",x"48"),
  1704 => (x"c2",x"87",x"ca",x"ff"),
  1705 => (x"6c",x"97",x"49",x"a5"),
  1706 => (x"4b",x"a3",x"71",x"4b"),
  1707 => (x"97",x"4b",x"6b",x"97"),
  1708 => (x"48",x"6e",x"7e",x"6c"),
  1709 => (x"a6",x"c8",x"80",x"c1"),
  1710 => (x"cc",x"98",x"c7",x"58"),
  1711 => (x"97",x"70",x"58",x"a6"),
  1712 => (x"87",x"e1",x"fe",x"7c"),
  1713 => (x"8e",x"f4",x"48",x"73"),
  1714 => (x"4c",x"26",x"4d",x"26"),
  1715 => (x"4f",x"26",x"4b",x"26"),
  1716 => (x"5c",x"5b",x"5e",x"0e"),
  1717 => (x"71",x"86",x"f4",x"0e"),
  1718 => (x"4a",x"66",x"d8",x"4c"),
  1719 => (x"c2",x"9a",x"ff",x"c3"),
  1720 => (x"6c",x"97",x"4b",x"a4"),
  1721 => (x"49",x"a1",x"73",x"49"),
  1722 => (x"6c",x"97",x"51",x"72"),
  1723 => (x"c1",x"48",x"6e",x"7e"),
  1724 => (x"58",x"a6",x"c8",x"80"),
  1725 => (x"a6",x"cc",x"98",x"c7"),
  1726 => (x"f4",x"54",x"70",x"58"),
  1727 => (x"87",x"ca",x"ff",x"8e"),
  1728 => (x"e8",x"fd",x"1e",x"1e"),
  1729 => (x"4a",x"bf",x"e0",x"87"),
  1730 => (x"c0",x"e0",x"c0",x"49"),
  1731 => (x"87",x"cb",x"02",x"99"),
  1732 => (x"f7",x"c2",x"1e",x"72"),
  1733 => (x"f7",x"fe",x"49",x"d2"),
  1734 => (x"fc",x"86",x"c4",x"87"),
  1735 => (x"7e",x"70",x"87",x"fd"),
  1736 => (x"26",x"87",x"c2",x"fd"),
  1737 => (x"c2",x"1e",x"4f",x"26"),
  1738 => (x"fd",x"49",x"d2",x"f7"),
  1739 => (x"ec",x"c1",x"87",x"c7"),
  1740 => (x"da",x"fc",x"49",x"c0"),
  1741 => (x"87",x"c7",x"c4",x"87"),
  1742 => (x"ff",x"1e",x"4f",x"26"),
  1743 => (x"e1",x"c8",x"48",x"d0"),
  1744 => (x"48",x"d4",x"ff",x"78"),
  1745 => (x"66",x"c4",x"78",x"c5"),
  1746 => (x"c3",x"87",x"c3",x"02"),
  1747 => (x"66",x"c8",x"78",x"e0"),
  1748 => (x"ff",x"87",x"c6",x"02"),
  1749 => (x"f0",x"c3",x"48",x"d4"),
  1750 => (x"48",x"d4",x"ff",x"78"),
  1751 => (x"d0",x"ff",x"78",x"71"),
  1752 => (x"78",x"e1",x"c8",x"48"),
  1753 => (x"26",x"78",x"e0",x"c0"),
  1754 => (x"5b",x"5e",x"0e",x"4f"),
  1755 => (x"4c",x"71",x"0e",x"5c"),
  1756 => (x"49",x"d2",x"f7",x"c2"),
  1757 => (x"70",x"87",x"c6",x"fc"),
  1758 => (x"aa",x"b7",x"c0",x"4a"),
  1759 => (x"87",x"e2",x"c2",x"04"),
  1760 => (x"05",x"aa",x"f0",x"c3"),
  1761 => (x"f0",x"c1",x"87",x"c9"),
  1762 => (x"78",x"c1",x"48",x"ee"),
  1763 => (x"c3",x"87",x"c3",x"c2"),
  1764 => (x"c9",x"05",x"aa",x"e0"),
  1765 => (x"f2",x"f0",x"c1",x"87"),
  1766 => (x"c1",x"78",x"c1",x"48"),
  1767 => (x"f0",x"c1",x"87",x"f4"),
  1768 => (x"c6",x"02",x"bf",x"f2"),
  1769 => (x"a2",x"c0",x"c2",x"87"),
  1770 => (x"72",x"87",x"c2",x"4b"),
  1771 => (x"05",x"9c",x"74",x"4b"),
  1772 => (x"f0",x"c1",x"87",x"d1"),
  1773 => (x"c1",x"1e",x"bf",x"ee"),
  1774 => (x"1e",x"bf",x"f2",x"f0"),
  1775 => (x"f9",x"fd",x"49",x"72"),
  1776 => (x"c1",x"86",x"c8",x"87"),
  1777 => (x"02",x"bf",x"ee",x"f0"),
  1778 => (x"73",x"87",x"e0",x"c0"),
  1779 => (x"29",x"b7",x"c4",x"49"),
  1780 => (x"ce",x"f2",x"c1",x"91"),
  1781 => (x"cf",x"4a",x"73",x"81"),
  1782 => (x"c1",x"92",x"c2",x"9a"),
  1783 => (x"70",x"30",x"72",x"48"),
  1784 => (x"72",x"ba",x"ff",x"4a"),
  1785 => (x"70",x"98",x"69",x"48"),
  1786 => (x"73",x"87",x"db",x"79"),
  1787 => (x"29",x"b7",x"c4",x"49"),
  1788 => (x"ce",x"f2",x"c1",x"91"),
  1789 => (x"cf",x"4a",x"73",x"81"),
  1790 => (x"c3",x"92",x"c2",x"9a"),
  1791 => (x"70",x"30",x"72",x"48"),
  1792 => (x"b0",x"69",x"48",x"4a"),
  1793 => (x"f0",x"c1",x"79",x"70"),
  1794 => (x"78",x"c0",x"48",x"f2"),
  1795 => (x"48",x"ee",x"f0",x"c1"),
  1796 => (x"f7",x"c2",x"78",x"c0"),
  1797 => (x"e4",x"f9",x"49",x"d2"),
  1798 => (x"c0",x"4a",x"70",x"87"),
  1799 => (x"fd",x"03",x"aa",x"b7"),
  1800 => (x"48",x"c0",x"87",x"de"),
  1801 => (x"4d",x"26",x"87",x"c2"),
  1802 => (x"4b",x"26",x"4c",x"26"),
  1803 => (x"00",x"00",x"4f",x"26"),
  1804 => (x"00",x"00",x"00",x"00"),
  1805 => (x"71",x"1e",x"00",x"00"),
  1806 => (x"ec",x"fc",x"49",x"4a"),
  1807 => (x"1e",x"4f",x"26",x"87"),
  1808 => (x"49",x"72",x"4a",x"c0"),
  1809 => (x"f2",x"c1",x"91",x"c4"),
  1810 => (x"79",x"c0",x"81",x"ce"),
  1811 => (x"b7",x"d0",x"82",x"c1"),
  1812 => (x"87",x"ee",x"04",x"aa"),
  1813 => (x"5e",x"0e",x"4f",x"26"),
  1814 => (x"0e",x"5d",x"5c",x"5b"),
  1815 => (x"cc",x"f8",x"4d",x"71"),
  1816 => (x"c4",x"4a",x"75",x"87"),
  1817 => (x"c1",x"92",x"2a",x"b7"),
  1818 => (x"75",x"82",x"ce",x"f2"),
  1819 => (x"c2",x"9c",x"cf",x"4c"),
  1820 => (x"4b",x"49",x"6a",x"94"),
  1821 => (x"9b",x"c3",x"2b",x"74"),
  1822 => (x"30",x"74",x"48",x"c2"),
  1823 => (x"bc",x"ff",x"4c",x"70"),
  1824 => (x"98",x"71",x"48",x"74"),
  1825 => (x"dc",x"f7",x"7a",x"70"),
  1826 => (x"fe",x"48",x"73",x"87"),
  1827 => (x"00",x"00",x"87",x"d8"),
  1828 => (x"00",x"00",x"00",x"00"),
  1829 => (x"00",x"00",x"00",x"00"),
  1830 => (x"00",x"00",x"00",x"00"),
  1831 => (x"00",x"00",x"00",x"00"),
  1832 => (x"00",x"00",x"00",x"00"),
  1833 => (x"00",x"00",x"00",x"00"),
  1834 => (x"00",x"00",x"00",x"00"),
  1835 => (x"00",x"00",x"00",x"00"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"00",x"00",x"00",x"00"),
  1838 => (x"00",x"00",x"00",x"00"),
  1839 => (x"00",x"00",x"00",x"00"),
  1840 => (x"00",x"00",x"00",x"00"),
  1841 => (x"00",x"00",x"00",x"00"),
  1842 => (x"00",x"00",x"00",x"00"),
  1843 => (x"ff",x"1e",x"00",x"00"),
  1844 => (x"e1",x"c8",x"48",x"d0"),
  1845 => (x"ff",x"48",x"71",x"78"),
  1846 => (x"c4",x"78",x"08",x"d4"),
  1847 => (x"d4",x"ff",x"48",x"66"),
  1848 => (x"4f",x"26",x"78",x"08"),
  1849 => (x"c4",x"4a",x"71",x"1e"),
  1850 => (x"72",x"1e",x"49",x"66"),
  1851 => (x"87",x"de",x"ff",x"49"),
  1852 => (x"c0",x"48",x"d0",x"ff"),
  1853 => (x"26",x"26",x"78",x"e0"),
  1854 => (x"1e",x"73",x"1e",x"4f"),
  1855 => (x"66",x"c8",x"4b",x"71"),
  1856 => (x"4a",x"73",x"1e",x"49"),
  1857 => (x"49",x"a2",x"e0",x"c1"),
  1858 => (x"26",x"87",x"d9",x"ff"),
  1859 => (x"4d",x"26",x"87",x"c4"),
  1860 => (x"4b",x"26",x"4c",x"26"),
  1861 => (x"73",x"1e",x"4f",x"26"),
  1862 => (x"4b",x"4a",x"71",x"1e"),
  1863 => (x"03",x"ab",x"b7",x"c2"),
  1864 => (x"49",x"a3",x"87",x"c8"),
  1865 => (x"9a",x"ff",x"c3",x"4a"),
  1866 => (x"a3",x"ce",x"87",x"c7"),
  1867 => (x"ff",x"c3",x"4a",x"49"),
  1868 => (x"49",x"66",x"c8",x"9a"),
  1869 => (x"fe",x"49",x"72",x"1e"),
  1870 => (x"ff",x"26",x"87",x"ea"),
  1871 => (x"ff",x"1e",x"87",x"d4"),
  1872 => (x"ff",x"c3",x"4a",x"d4"),
  1873 => (x"48",x"d0",x"ff",x"7a"),
  1874 => (x"de",x"78",x"e1",x"c0"),
  1875 => (x"dc",x"f7",x"c2",x"7a"),
  1876 => (x"48",x"49",x"7a",x"bf"),
  1877 => (x"7a",x"70",x"28",x"c8"),
  1878 => (x"28",x"d0",x"48",x"71"),
  1879 => (x"48",x"71",x"7a",x"70"),
  1880 => (x"7a",x"70",x"28",x"d8"),
  1881 => (x"c0",x"48",x"d0",x"ff"),
  1882 => (x"4f",x"26",x"78",x"e0"),
  1883 => (x"5c",x"5b",x"5e",x"0e"),
  1884 => (x"4c",x"71",x"0e",x"5d"),
  1885 => (x"bf",x"dc",x"f7",x"c2"),
  1886 => (x"2b",x"74",x"4b",x"4d"),
  1887 => (x"c1",x"9b",x"66",x"d0"),
  1888 => (x"ab",x"66",x"d4",x"83"),
  1889 => (x"c0",x"87",x"c2",x"04"),
  1890 => (x"d0",x"4a",x"74",x"4b"),
  1891 => (x"31",x"72",x"49",x"66"),
  1892 => (x"99",x"75",x"b9",x"ff"),
  1893 => (x"30",x"72",x"48",x"73"),
  1894 => (x"71",x"48",x"4a",x"70"),
  1895 => (x"e0",x"f7",x"c2",x"b0"),
  1896 => (x"87",x"da",x"fe",x"58"),
  1897 => (x"4c",x"26",x"4d",x"26"),
  1898 => (x"4f",x"26",x"4b",x"26"),
  1899 => (x"5c",x"5b",x"5e",x"0e"),
  1900 => (x"71",x"1e",x"0e",x"5d"),
  1901 => (x"e0",x"f7",x"c2",x"4c"),
  1902 => (x"c0",x"4a",x"c0",x"4b"),
  1903 => (x"cc",x"fe",x"49",x"f4"),
  1904 => (x"1e",x"74",x"87",x"c3"),
  1905 => (x"49",x"e0",x"f7",x"c2"),
  1906 => (x"87",x"c6",x"e7",x"fe"),
  1907 => (x"49",x"70",x"86",x"c4"),
  1908 => (x"ea",x"c0",x"02",x"99"),
  1909 => (x"a6",x"1e",x"c4",x"87"),
  1910 => (x"f7",x"c2",x"1e",x"4d"),
  1911 => (x"ee",x"fe",x"49",x"e0"),
  1912 => (x"86",x"c8",x"87",x"d9"),
  1913 => (x"d6",x"02",x"98",x"70"),
  1914 => (x"c1",x"4a",x"75",x"87"),
  1915 => (x"c4",x"49",x"f5",x"f8"),
  1916 => (x"f5",x"c9",x"fe",x"4b"),
  1917 => (x"02",x"98",x"70",x"87"),
  1918 => (x"48",x"c0",x"87",x"ca"),
  1919 => (x"c0",x"87",x"ed",x"c0"),
  1920 => (x"87",x"e8",x"c0",x"48"),
  1921 => (x"c1",x"87",x"f3",x"c0"),
  1922 => (x"98",x"70",x"87",x"c4"),
  1923 => (x"c0",x"87",x"c8",x"02"),
  1924 => (x"98",x"70",x"87",x"fc"),
  1925 => (x"c2",x"87",x"f8",x"05"),
  1926 => (x"02",x"bf",x"c0",x"f8"),
  1927 => (x"f7",x"c2",x"87",x"cc"),
  1928 => (x"f8",x"c2",x"48",x"dc"),
  1929 => (x"fc",x"78",x"bf",x"c0"),
  1930 => (x"48",x"c1",x"87",x"d4"),
  1931 => (x"26",x"4d",x"26",x"26"),
  1932 => (x"26",x"4b",x"26",x"4c"),
  1933 => (x"52",x"41",x"5b",x"4f"),
  1934 => (x"c0",x"1e",x"00",x"43"),
  1935 => (x"e0",x"f7",x"c2",x"1e"),
  1936 => (x"cf",x"eb",x"fe",x"49"),
  1937 => (x"f8",x"f7",x"c2",x"87"),
  1938 => (x"26",x"78",x"c0",x"48"),
  1939 => (x"5e",x"0e",x"4f",x"26"),
  1940 => (x"0e",x"5d",x"5c",x"5b"),
  1941 => (x"a6",x"c4",x"86",x"f4"),
  1942 => (x"c2",x"78",x"c0",x"48"),
  1943 => (x"48",x"bf",x"f8",x"f7"),
  1944 => (x"03",x"a8",x"b7",x"c3"),
  1945 => (x"f7",x"c2",x"87",x"d1"),
  1946 => (x"c1",x"48",x"bf",x"f8"),
  1947 => (x"fc",x"f7",x"c2",x"80"),
  1948 => (x"48",x"fb",x"c0",x"58"),
  1949 => (x"c2",x"87",x"e2",x"c6"),
  1950 => (x"fe",x"49",x"e0",x"f7"),
  1951 => (x"70",x"87",x"d0",x"f0"),
  1952 => (x"f8",x"f7",x"c2",x"4c"),
  1953 => (x"8a",x"c3",x"4a",x"bf"),
  1954 => (x"c1",x"87",x"d8",x"02"),
  1955 => (x"cb",x"c5",x"02",x"8a"),
  1956 => (x"c2",x"02",x"8a",x"87"),
  1957 => (x"02",x"8a",x"87",x"f6"),
  1958 => (x"8a",x"87",x"cd",x"c1"),
  1959 => (x"87",x"e2",x"c3",x"02"),
  1960 => (x"c0",x"87",x"e1",x"c5"),
  1961 => (x"c4",x"4a",x"75",x"4d"),
  1962 => (x"f7",x"c0",x"c2",x"92"),
  1963 => (x"f4",x"f7",x"c2",x"82"),
  1964 => (x"70",x"80",x"75",x"48"),
  1965 => (x"bf",x"97",x"6e",x"7e"),
  1966 => (x"6e",x"4b",x"49",x"4b"),
  1967 => (x"50",x"a3",x"c1",x"48"),
  1968 => (x"48",x"11",x"81",x"6a"),
  1969 => (x"70",x"58",x"a6",x"cc"),
  1970 => (x"87",x"c4",x"02",x"ac"),
  1971 => (x"50",x"c0",x"48",x"6e"),
  1972 => (x"c7",x"05",x"66",x"c8"),
  1973 => (x"f8",x"f7",x"c2",x"87"),
  1974 => (x"78",x"a5",x"c4",x"48"),
  1975 => (x"b7",x"c4",x"85",x"c1"),
  1976 => (x"c0",x"ff",x"04",x"ad"),
  1977 => (x"87",x"dc",x"c4",x"87"),
  1978 => (x"bf",x"c4",x"f8",x"c2"),
  1979 => (x"a8",x"b7",x"c8",x"48"),
  1980 => (x"ca",x"87",x"d1",x"01"),
  1981 => (x"87",x"cc",x"02",x"ac"),
  1982 => (x"c7",x"02",x"ac",x"cd"),
  1983 => (x"ac",x"b7",x"c0",x"87"),
  1984 => (x"87",x"f3",x"c0",x"03"),
  1985 => (x"bf",x"c4",x"f8",x"c2"),
  1986 => (x"ab",x"b7",x"c8",x"4b"),
  1987 => (x"c2",x"87",x"d2",x"03"),
  1988 => (x"73",x"49",x"c8",x"f8"),
  1989 => (x"51",x"e0",x"c0",x"81"),
  1990 => (x"b7",x"c8",x"83",x"c1"),
  1991 => (x"ee",x"ff",x"04",x"ab"),
  1992 => (x"d0",x"f8",x"c2",x"87"),
  1993 => (x"50",x"d2",x"c1",x"48"),
  1994 => (x"c1",x"50",x"cf",x"c1"),
  1995 => (x"50",x"c0",x"50",x"cd"),
  1996 => (x"78",x"c3",x"80",x"e4"),
  1997 => (x"c2",x"87",x"cd",x"c3"),
  1998 => (x"49",x"bf",x"c4",x"f8"),
  1999 => (x"c2",x"80",x"c1",x"48"),
  2000 => (x"48",x"58",x"c8",x"f8"),
  2001 => (x"74",x"81",x"a0",x"c4"),
  2002 => (x"87",x"f8",x"c2",x"51"),
  2003 => (x"ac",x"b7",x"f0",x"c0"),
  2004 => (x"c0",x"87",x"da",x"04"),
  2005 => (x"01",x"ac",x"b7",x"f9"),
  2006 => (x"f7",x"c2",x"87",x"d3"),
  2007 => (x"ca",x"49",x"bf",x"fc"),
  2008 => (x"c0",x"4a",x"74",x"91"),
  2009 => (x"f7",x"c2",x"8a",x"f0"),
  2010 => (x"a1",x"72",x"48",x"fc"),
  2011 => (x"02",x"ac",x"ca",x"78"),
  2012 => (x"cd",x"87",x"c6",x"c0"),
  2013 => (x"cb",x"c2",x"05",x"ac"),
  2014 => (x"f8",x"f7",x"c2",x"87"),
  2015 => (x"c2",x"78",x"c3",x"48"),
  2016 => (x"f0",x"c0",x"87",x"c2"),
  2017 => (x"db",x"04",x"ac",x"b7"),
  2018 => (x"b7",x"f9",x"c0",x"87"),
  2019 => (x"d3",x"c0",x"01",x"ac"),
  2020 => (x"c0",x"f8",x"c2",x"87"),
  2021 => (x"91",x"d0",x"49",x"bf"),
  2022 => (x"f0",x"c0",x"4a",x"74"),
  2023 => (x"c0",x"f8",x"c2",x"8a"),
  2024 => (x"78",x"a1",x"72",x"48"),
  2025 => (x"ac",x"b7",x"c1",x"c1"),
  2026 => (x"87",x"db",x"c0",x"04"),
  2027 => (x"ac",x"b7",x"c6",x"c1"),
  2028 => (x"87",x"d3",x"c0",x"01"),
  2029 => (x"bf",x"c0",x"f8",x"c2"),
  2030 => (x"74",x"91",x"d0",x"49"),
  2031 => (x"8a",x"f7",x"c0",x"4a"),
  2032 => (x"48",x"c0",x"f8",x"c2"),
  2033 => (x"ca",x"78",x"a1",x"72"),
  2034 => (x"c6",x"c0",x"02",x"ac"),
  2035 => (x"05",x"ac",x"cd",x"87"),
  2036 => (x"c2",x"87",x"f1",x"c0"),
  2037 => (x"c3",x"48",x"f8",x"f7"),
  2038 => (x"87",x"e8",x"c0",x"78"),
  2039 => (x"05",x"ac",x"e2",x"c0"),
  2040 => (x"c4",x"87",x"c9",x"c0"),
  2041 => (x"fb",x"c0",x"48",x"a6"),
  2042 => (x"87",x"d8",x"c0",x"78"),
  2043 => (x"c0",x"02",x"ac",x"ca"),
  2044 => (x"ac",x"cd",x"87",x"c6"),
  2045 => (x"87",x"c9",x"c0",x"05"),
  2046 => (x"48",x"f8",x"f7",x"c2"),
  2047 => (x"c3",x"c0",x"78",x"c3"),
  2048 => (x"5c",x"a6",x"c8",x"87"),
  2049 => (x"03",x"ac",x"b7",x"c0"),
  2050 => (x"48",x"87",x"c4",x"c0"),
  2051 => (x"c4",x"87",x"ca",x"c0"),
  2052 => (x"c6",x"f9",x"02",x"66"),
  2053 => (x"ff",x"c3",x"48",x"87"),
  2054 => (x"f8",x"8e",x"f4",x"99"),
  2055 => (x"4f",x"43",x"87",x"cf"),
  2056 => (x"00",x"3d",x"46",x"4e"),
  2057 => (x"00",x"44",x"4f",x"4d"),
  2058 => (x"45",x"4d",x"41",x"4e"),
  2059 => (x"46",x"45",x"44",x"00"),
  2060 => (x"54",x"4c",x"55",x"41"),
  2061 => (x"1e",x"00",x"30",x"3d"),
  2062 => (x"24",x"00",x"00",x"20"),
  2063 => (x"28",x"00",x"00",x"20"),
  2064 => (x"2d",x"00",x"00",x"20"),
  2065 => (x"1e",x"00",x"00",x"20"),
  2066 => (x"c8",x"48",x"d0",x"ff"),
  2067 => (x"48",x"71",x"78",x"c9"),
  2068 => (x"78",x"08",x"d4",x"ff"),
  2069 => (x"71",x"1e",x"4f",x"26"),
  2070 => (x"87",x"eb",x"49",x"4a"),
  2071 => (x"c8",x"48",x"d0",x"ff"),
  2072 => (x"1e",x"4f",x"26",x"78"),
  2073 => (x"4b",x"71",x"1e",x"73"),
  2074 => (x"bf",x"e0",x"f8",x"c2"),
  2075 => (x"c2",x"87",x"c3",x"02"),
  2076 => (x"d0",x"ff",x"87",x"eb"),
  2077 => (x"78",x"c9",x"c8",x"48"),
  2078 => (x"e0",x"c0",x"49",x"73"),
  2079 => (x"48",x"d4",x"ff",x"b1"),
  2080 => (x"f8",x"c2",x"78",x"71"),
  2081 => (x"78",x"c0",x"48",x"d4"),
  2082 => (x"c5",x"02",x"66",x"c8"),
  2083 => (x"49",x"ff",x"c3",x"87"),
  2084 => (x"49",x"c0",x"87",x"c2"),
  2085 => (x"59",x"dc",x"f8",x"c2"),
  2086 => (x"c6",x"02",x"66",x"cc"),
  2087 => (x"d5",x"d5",x"c5",x"87"),
  2088 => (x"cf",x"87",x"c4",x"4a"),
  2089 => (x"c2",x"4a",x"ff",x"ff"),
  2090 => (x"c2",x"5a",x"e0",x"f8"),
  2091 => (x"c1",x"48",x"e0",x"f8"),
  2092 => (x"26",x"87",x"c4",x"78"),
  2093 => (x"26",x"4c",x"26",x"4d"),
  2094 => (x"0e",x"4f",x"26",x"4b"),
  2095 => (x"5d",x"5c",x"5b",x"5e"),
  2096 => (x"c2",x"4a",x"71",x"0e"),
  2097 => (x"4c",x"bf",x"dc",x"f8"),
  2098 => (x"cb",x"02",x"9a",x"72"),
  2099 => (x"91",x"c8",x"49",x"87"),
  2100 => (x"4b",x"d9",x"c1",x"c2"),
  2101 => (x"87",x"c4",x"83",x"71"),
  2102 => (x"4b",x"d9",x"c5",x"c2"),
  2103 => (x"49",x"13",x"4d",x"c0"),
  2104 => (x"f8",x"c2",x"99",x"74"),
  2105 => (x"ff",x"b9",x"bf",x"d8"),
  2106 => (x"78",x"71",x"48",x"d4"),
  2107 => (x"85",x"2c",x"b7",x"c1"),
  2108 => (x"04",x"ad",x"b7",x"c8"),
  2109 => (x"f8",x"c2",x"87",x"e8"),
  2110 => (x"c8",x"48",x"bf",x"d4"),
  2111 => (x"d8",x"f8",x"c2",x"80"),
  2112 => (x"87",x"ef",x"fe",x"58"),
  2113 => (x"71",x"1e",x"73",x"1e"),
  2114 => (x"9a",x"4a",x"13",x"4b"),
  2115 => (x"72",x"87",x"cb",x"02"),
  2116 => (x"87",x"e7",x"fe",x"49"),
  2117 => (x"05",x"9a",x"4a",x"13"),
  2118 => (x"da",x"fe",x"87",x"f5"),
  2119 => (x"f8",x"c2",x"1e",x"87"),
  2120 => (x"c2",x"49",x"bf",x"d4"),
  2121 => (x"c1",x"48",x"d4",x"f8"),
  2122 => (x"c0",x"c4",x"78",x"a1"),
  2123 => (x"db",x"03",x"a9",x"b7"),
  2124 => (x"48",x"d4",x"ff",x"87"),
  2125 => (x"bf",x"d8",x"f8",x"c2"),
  2126 => (x"d4",x"f8",x"c2",x"78"),
  2127 => (x"f8",x"c2",x"49",x"bf"),
  2128 => (x"a1",x"c1",x"48",x"d4"),
  2129 => (x"b7",x"c0",x"c4",x"78"),
  2130 => (x"87",x"e5",x"04",x"a9"),
  2131 => (x"c8",x"48",x"d0",x"ff"),
  2132 => (x"e0",x"f8",x"c2",x"78"),
  2133 => (x"26",x"78",x"c0",x"48"),
  2134 => (x"00",x"00",x"00",x"4f"),
  2135 => (x"00",x"00",x"00",x"00"),
  2136 => (x"00",x"00",x"00",x"00"),
  2137 => (x"00",x"00",x"5f",x"5f"),
  2138 => (x"03",x"03",x"00",x"00"),
  2139 => (x"00",x"03",x"03",x"00"),
  2140 => (x"7f",x"7f",x"14",x"00"),
  2141 => (x"14",x"7f",x"7f",x"14"),
  2142 => (x"2e",x"24",x"00",x"00"),
  2143 => (x"12",x"3a",x"6b",x"6b"),
  2144 => (x"36",x"6a",x"4c",x"00"),
  2145 => (x"32",x"56",x"6c",x"18"),
  2146 => (x"4f",x"7e",x"30",x"00"),
  2147 => (x"68",x"3a",x"77",x"59"),
  2148 => (x"04",x"00",x"00",x"40"),
  2149 => (x"00",x"00",x"03",x"07"),
  2150 => (x"1c",x"00",x"00",x"00"),
  2151 => (x"00",x"41",x"63",x"3e"),
  2152 => (x"41",x"00",x"00",x"00"),
  2153 => (x"00",x"1c",x"3e",x"63"),
  2154 => (x"3e",x"2a",x"08",x"00"),
  2155 => (x"2a",x"3e",x"1c",x"1c"),
  2156 => (x"08",x"08",x"00",x"08"),
  2157 => (x"08",x"08",x"3e",x"3e"),
  2158 => (x"80",x"00",x"00",x"00"),
  2159 => (x"00",x"00",x"60",x"e0"),
  2160 => (x"08",x"08",x"00",x"00"),
  2161 => (x"08",x"08",x"08",x"08"),
  2162 => (x"00",x"00",x"00",x"00"),
  2163 => (x"00",x"00",x"60",x"60"),
  2164 => (x"30",x"60",x"40",x"00"),
  2165 => (x"03",x"06",x"0c",x"18"),
  2166 => (x"7f",x"3e",x"00",x"01"),
  2167 => (x"3e",x"7f",x"4d",x"59"),
  2168 => (x"06",x"04",x"00",x"00"),
  2169 => (x"00",x"00",x"7f",x"7f"),
  2170 => (x"63",x"42",x"00",x"00"),
  2171 => (x"46",x"4f",x"59",x"71"),
  2172 => (x"63",x"22",x"00",x"00"),
  2173 => (x"36",x"7f",x"49",x"49"),
  2174 => (x"16",x"1c",x"18",x"00"),
  2175 => (x"10",x"7f",x"7f",x"13"),
  2176 => (x"67",x"27",x"00",x"00"),
  2177 => (x"39",x"7d",x"45",x"45"),
  2178 => (x"7e",x"3c",x"00",x"00"),
  2179 => (x"30",x"79",x"49",x"4b"),
  2180 => (x"01",x"01",x"00",x"00"),
  2181 => (x"07",x"0f",x"79",x"71"),
  2182 => (x"7f",x"36",x"00",x"00"),
  2183 => (x"36",x"7f",x"49",x"49"),
  2184 => (x"4f",x"06",x"00",x"00"),
  2185 => (x"1e",x"3f",x"69",x"49"),
  2186 => (x"00",x"00",x"00",x"00"),
  2187 => (x"00",x"00",x"66",x"66"),
  2188 => (x"80",x"00",x"00",x"00"),
  2189 => (x"00",x"00",x"66",x"e6"),
  2190 => (x"08",x"08",x"00",x"00"),
  2191 => (x"22",x"22",x"14",x"14"),
  2192 => (x"14",x"14",x"00",x"00"),
  2193 => (x"14",x"14",x"14",x"14"),
  2194 => (x"22",x"22",x"00",x"00"),
  2195 => (x"08",x"08",x"14",x"14"),
  2196 => (x"03",x"02",x"00",x"00"),
  2197 => (x"06",x"0f",x"59",x"51"),
  2198 => (x"41",x"7f",x"3e",x"00"),
  2199 => (x"1e",x"1f",x"55",x"5d"),
  2200 => (x"7f",x"7e",x"00",x"00"),
  2201 => (x"7e",x"7f",x"09",x"09"),
  2202 => (x"7f",x"7f",x"00",x"00"),
  2203 => (x"36",x"7f",x"49",x"49"),
  2204 => (x"3e",x"1c",x"00",x"00"),
  2205 => (x"41",x"41",x"41",x"63"),
  2206 => (x"7f",x"7f",x"00",x"00"),
  2207 => (x"1c",x"3e",x"63",x"41"),
  2208 => (x"7f",x"7f",x"00",x"00"),
  2209 => (x"41",x"41",x"49",x"49"),
  2210 => (x"7f",x"7f",x"00",x"00"),
  2211 => (x"01",x"01",x"09",x"09"),
  2212 => (x"7f",x"3e",x"00",x"00"),
  2213 => (x"7a",x"7b",x"49",x"41"),
  2214 => (x"7f",x"7f",x"00",x"00"),
  2215 => (x"7f",x"7f",x"08",x"08"),
  2216 => (x"41",x"00",x"00",x"00"),
  2217 => (x"00",x"41",x"7f",x"7f"),
  2218 => (x"60",x"20",x"00",x"00"),
  2219 => (x"3f",x"7f",x"40",x"40"),
  2220 => (x"08",x"7f",x"7f",x"00"),
  2221 => (x"41",x"63",x"36",x"1c"),
  2222 => (x"7f",x"7f",x"00",x"00"),
  2223 => (x"40",x"40",x"40",x"40"),
  2224 => (x"06",x"7f",x"7f",x"00"),
  2225 => (x"7f",x"7f",x"06",x"0c"),
  2226 => (x"06",x"7f",x"7f",x"00"),
  2227 => (x"7f",x"7f",x"18",x"0c"),
  2228 => (x"7f",x"3e",x"00",x"00"),
  2229 => (x"3e",x"7f",x"41",x"41"),
  2230 => (x"7f",x"7f",x"00",x"00"),
  2231 => (x"06",x"0f",x"09",x"09"),
  2232 => (x"41",x"7f",x"3e",x"00"),
  2233 => (x"40",x"7e",x"7f",x"61"),
  2234 => (x"7f",x"7f",x"00",x"00"),
  2235 => (x"66",x"7f",x"19",x"09"),
  2236 => (x"6f",x"26",x"00",x"00"),
  2237 => (x"32",x"7b",x"59",x"4d"),
  2238 => (x"01",x"01",x"00",x"00"),
  2239 => (x"01",x"01",x"7f",x"7f"),
  2240 => (x"7f",x"3f",x"00",x"00"),
  2241 => (x"3f",x"7f",x"40",x"40"),
  2242 => (x"3f",x"0f",x"00",x"00"),
  2243 => (x"0f",x"3f",x"70",x"70"),
  2244 => (x"30",x"7f",x"7f",x"00"),
  2245 => (x"7f",x"7f",x"30",x"18"),
  2246 => (x"36",x"63",x"41",x"00"),
  2247 => (x"63",x"36",x"1c",x"1c"),
  2248 => (x"06",x"03",x"01",x"41"),
  2249 => (x"03",x"06",x"7c",x"7c"),
  2250 => (x"59",x"71",x"61",x"01"),
  2251 => (x"41",x"43",x"47",x"4d"),
  2252 => (x"7f",x"00",x"00",x"00"),
  2253 => (x"00",x"41",x"41",x"7f"),
  2254 => (x"06",x"03",x"01",x"00"),
  2255 => (x"60",x"30",x"18",x"0c"),
  2256 => (x"41",x"00",x"00",x"40"),
  2257 => (x"00",x"7f",x"7f",x"41"),
  2258 => (x"06",x"0c",x"08",x"00"),
  2259 => (x"08",x"0c",x"06",x"03"),
  2260 => (x"80",x"80",x"80",x"00"),
  2261 => (x"80",x"80",x"80",x"80"),
  2262 => (x"00",x"00",x"00",x"00"),
  2263 => (x"00",x"04",x"07",x"03"),
  2264 => (x"74",x"20",x"00",x"00"),
  2265 => (x"78",x"7c",x"54",x"54"),
  2266 => (x"7f",x"7f",x"00",x"00"),
  2267 => (x"38",x"7c",x"44",x"44"),
  2268 => (x"7c",x"38",x"00",x"00"),
  2269 => (x"00",x"44",x"44",x"44"),
  2270 => (x"7c",x"38",x"00",x"00"),
  2271 => (x"7f",x"7f",x"44",x"44"),
  2272 => (x"7c",x"38",x"00",x"00"),
  2273 => (x"18",x"5c",x"54",x"54"),
  2274 => (x"7e",x"04",x"00",x"00"),
  2275 => (x"00",x"05",x"05",x"7f"),
  2276 => (x"bc",x"18",x"00",x"00"),
  2277 => (x"7c",x"fc",x"a4",x"a4"),
  2278 => (x"7f",x"7f",x"00",x"00"),
  2279 => (x"78",x"7c",x"04",x"04"),
  2280 => (x"00",x"00",x"00",x"00"),
  2281 => (x"00",x"40",x"7d",x"3d"),
  2282 => (x"80",x"80",x"00",x"00"),
  2283 => (x"00",x"7d",x"fd",x"80"),
  2284 => (x"7f",x"7f",x"00",x"00"),
  2285 => (x"44",x"6c",x"38",x"10"),
  2286 => (x"00",x"00",x"00",x"00"),
  2287 => (x"00",x"40",x"7f",x"3f"),
  2288 => (x"0c",x"7c",x"7c",x"00"),
  2289 => (x"78",x"7c",x"0c",x"18"),
  2290 => (x"7c",x"7c",x"00",x"00"),
  2291 => (x"78",x"7c",x"04",x"04"),
  2292 => (x"7c",x"38",x"00",x"00"),
  2293 => (x"38",x"7c",x"44",x"44"),
  2294 => (x"fc",x"fc",x"00",x"00"),
  2295 => (x"18",x"3c",x"24",x"24"),
  2296 => (x"3c",x"18",x"00",x"00"),
  2297 => (x"fc",x"fc",x"24",x"24"),
  2298 => (x"7c",x"7c",x"00",x"00"),
  2299 => (x"08",x"0c",x"04",x"04"),
  2300 => (x"5c",x"48",x"00",x"00"),
  2301 => (x"20",x"74",x"54",x"54"),
  2302 => (x"3f",x"04",x"00",x"00"),
  2303 => (x"00",x"44",x"44",x"7f"),
  2304 => (x"7c",x"3c",x"00",x"00"),
  2305 => (x"7c",x"7c",x"40",x"40"),
  2306 => (x"3c",x"1c",x"00",x"00"),
  2307 => (x"1c",x"3c",x"60",x"60"),
  2308 => (x"60",x"7c",x"3c",x"00"),
  2309 => (x"3c",x"7c",x"60",x"30"),
  2310 => (x"38",x"6c",x"44",x"00"),
  2311 => (x"44",x"6c",x"38",x"10"),
  2312 => (x"bc",x"1c",x"00",x"00"),
  2313 => (x"1c",x"3c",x"60",x"e0"),
  2314 => (x"64",x"44",x"00",x"00"),
  2315 => (x"44",x"4c",x"5c",x"74"),
  2316 => (x"08",x"08",x"00",x"00"),
  2317 => (x"41",x"41",x"77",x"3e"),
  2318 => (x"00",x"00",x"00",x"00"),
  2319 => (x"00",x"00",x"7f",x"7f"),
  2320 => (x"41",x"41",x"00",x"00"),
  2321 => (x"08",x"08",x"3e",x"77"),
  2322 => (x"01",x"01",x"02",x"00"),
  2323 => (x"01",x"02",x"02",x"03"),
  2324 => (x"7f",x"7f",x"7f",x"00"),
  2325 => (x"7f",x"7f",x"7f",x"7f"),
  2326 => (x"1c",x"08",x"08",x"00"),
  2327 => (x"7f",x"3e",x"3e",x"1c"),
  2328 => (x"3e",x"7f",x"7f",x"7f"),
  2329 => (x"08",x"1c",x"1c",x"3e"),
  2330 => (x"18",x"10",x"00",x"08"),
  2331 => (x"10",x"18",x"7c",x"7c"),
  2332 => (x"30",x"10",x"00",x"00"),
  2333 => (x"10",x"30",x"7c",x"7c"),
  2334 => (x"60",x"30",x"10",x"00"),
  2335 => (x"06",x"1e",x"78",x"60"),
  2336 => (x"3c",x"66",x"42",x"00"),
  2337 => (x"42",x"66",x"3c",x"18"),
  2338 => (x"6a",x"38",x"78",x"00"),
  2339 => (x"38",x"6c",x"c6",x"c2"),
  2340 => (x"00",x"00",x"60",x"00"),
  2341 => (x"60",x"00",x"00",x"60"),
  2342 => (x"5b",x"5e",x"0e",x"00"),
  2343 => (x"1e",x"0e",x"5d",x"5c"),
  2344 => (x"f8",x"c2",x"4c",x"71"),
  2345 => (x"c0",x"4d",x"bf",x"f1"),
  2346 => (x"74",x"1e",x"c0",x"4b"),
  2347 => (x"87",x"c7",x"02",x"ab"),
  2348 => (x"c0",x"48",x"a6",x"c4"),
  2349 => (x"c4",x"87",x"c5",x"78"),
  2350 => (x"78",x"c1",x"48",x"a6"),
  2351 => (x"73",x"1e",x"66",x"c4"),
  2352 => (x"87",x"df",x"ee",x"49"),
  2353 => (x"e0",x"c0",x"86",x"c8"),
  2354 => (x"87",x"ef",x"ef",x"49"),
  2355 => (x"6a",x"4a",x"a5",x"c4"),
  2356 => (x"87",x"f0",x"f0",x"49"),
  2357 => (x"cb",x"87",x"c6",x"f1"),
  2358 => (x"c8",x"83",x"c1",x"85"),
  2359 => (x"ff",x"04",x"ab",x"b7"),
  2360 => (x"26",x"26",x"87",x"c7"),
  2361 => (x"26",x"4c",x"26",x"4d"),
  2362 => (x"1e",x"4f",x"26",x"4b"),
  2363 => (x"f8",x"c2",x"4a",x"71"),
  2364 => (x"f8",x"c2",x"5a",x"f5"),
  2365 => (x"78",x"c7",x"48",x"f5"),
  2366 => (x"87",x"dd",x"fe",x"49"),
  2367 => (x"73",x"1e",x"4f",x"26"),
  2368 => (x"c0",x"4a",x"71",x"1e"),
  2369 => (x"d3",x"03",x"aa",x"b7"),
  2370 => (x"de",x"e1",x"c2",x"87"),
  2371 => (x"87",x"c4",x"05",x"bf"),
  2372 => (x"87",x"c2",x"4b",x"c1"),
  2373 => (x"e1",x"c2",x"4b",x"c0"),
  2374 => (x"87",x"c4",x"5b",x"e2"),
  2375 => (x"5a",x"e2",x"e1",x"c2"),
  2376 => (x"bf",x"de",x"e1",x"c2"),
  2377 => (x"c1",x"9a",x"c1",x"4a"),
  2378 => (x"ec",x"49",x"a2",x"c0"),
  2379 => (x"48",x"fc",x"87",x"e8"),
  2380 => (x"bf",x"de",x"e1",x"c2"),
  2381 => (x"87",x"ef",x"fe",x"78"),
  2382 => (x"c4",x"4a",x"71",x"1e"),
  2383 => (x"49",x"72",x"1e",x"66"),
  2384 => (x"87",x"d2",x"df",x"ff"),
  2385 => (x"1e",x"4f",x"26",x"26"),
  2386 => (x"bf",x"de",x"e1",x"c2"),
  2387 => (x"e5",x"db",x"ff",x"49"),
  2388 => (x"e9",x"f8",x"c2",x"87"),
  2389 => (x"78",x"bf",x"e8",x"48"),
  2390 => (x"48",x"e5",x"f8",x"c2"),
  2391 => (x"c2",x"78",x"bf",x"ec"),
  2392 => (x"4a",x"bf",x"e9",x"f8"),
  2393 => (x"99",x"ff",x"c3",x"49"),
  2394 => (x"72",x"2a",x"b7",x"c8"),
  2395 => (x"c2",x"b0",x"71",x"48"),
  2396 => (x"26",x"58",x"f1",x"f8"),
  2397 => (x"5b",x"5e",x"0e",x"4f"),
  2398 => (x"71",x"0e",x"5d",x"5c"),
  2399 => (x"87",x"c7",x"ff",x"4b"),
  2400 => (x"48",x"e4",x"f8",x"c2"),
  2401 => (x"49",x"73",x"50",x"c0"),
  2402 => (x"87",x"ca",x"db",x"ff"),
  2403 => (x"c2",x"4c",x"49",x"70"),
  2404 => (x"49",x"ee",x"cb",x"9c"),
  2405 => (x"70",x"87",x"cf",x"cb"),
  2406 => (x"f8",x"c2",x"4d",x"49"),
  2407 => (x"05",x"bf",x"97",x"e4"),
  2408 => (x"d0",x"87",x"e4",x"c1"),
  2409 => (x"f8",x"c2",x"49",x"66"),
  2410 => (x"05",x"99",x"bf",x"ed"),
  2411 => (x"66",x"d4",x"87",x"d7"),
  2412 => (x"e5",x"f8",x"c2",x"49"),
  2413 => (x"cc",x"05",x"99",x"bf"),
  2414 => (x"ff",x"49",x"73",x"87"),
  2415 => (x"70",x"87",x"d7",x"da"),
  2416 => (x"c2",x"c1",x"02",x"98"),
  2417 => (x"fd",x"4c",x"c1",x"87"),
  2418 => (x"49",x"75",x"87",x"fd"),
  2419 => (x"70",x"87",x"e3",x"ca"),
  2420 => (x"87",x"c6",x"02",x"98"),
  2421 => (x"48",x"e4",x"f8",x"c2"),
  2422 => (x"f8",x"c2",x"50",x"c1"),
  2423 => (x"05",x"bf",x"97",x"e4"),
  2424 => (x"c2",x"87",x"e4",x"c0"),
  2425 => (x"49",x"bf",x"ed",x"f8"),
  2426 => (x"05",x"99",x"66",x"d0"),
  2427 => (x"c2",x"87",x"d6",x"ff"),
  2428 => (x"49",x"bf",x"e5",x"f8"),
  2429 => (x"05",x"99",x"66",x"d4"),
  2430 => (x"73",x"87",x"ca",x"ff"),
  2431 => (x"d5",x"d9",x"ff",x"49"),
  2432 => (x"05",x"98",x"70",x"87"),
  2433 => (x"74",x"87",x"fe",x"fe"),
  2434 => (x"87",x"d7",x"fb",x"48"),
  2435 => (x"5c",x"5b",x"5e",x"0e"),
  2436 => (x"86",x"f4",x"0e",x"5d"),
  2437 => (x"ec",x"4c",x"4d",x"c0"),
  2438 => (x"a6",x"c4",x"7e",x"bf"),
  2439 => (x"f1",x"f8",x"c2",x"48"),
  2440 => (x"1e",x"c1",x"78",x"bf"),
  2441 => (x"49",x"c7",x"1e",x"c0"),
  2442 => (x"c8",x"87",x"ca",x"fd"),
  2443 => (x"02",x"98",x"70",x"86"),
  2444 => (x"49",x"ff",x"87",x"ce"),
  2445 => (x"c1",x"87",x"c7",x"fb"),
  2446 => (x"d8",x"ff",x"49",x"da"),
  2447 => (x"4d",x"c1",x"87",x"d8"),
  2448 => (x"97",x"e4",x"f8",x"c2"),
  2449 => (x"87",x"c3",x"02",x"bf"),
  2450 => (x"c2",x"87",x"c0",x"c9"),
  2451 => (x"4b",x"bf",x"e9",x"f8"),
  2452 => (x"bf",x"de",x"e1",x"c2"),
  2453 => (x"87",x"eb",x"c0",x"05"),
  2454 => (x"ff",x"49",x"fd",x"c3"),
  2455 => (x"c3",x"87",x"f7",x"d7"),
  2456 => (x"d7",x"ff",x"49",x"fa"),
  2457 => (x"49",x"73",x"87",x"f0"),
  2458 => (x"71",x"99",x"ff",x"c3"),
  2459 => (x"fb",x"49",x"c0",x"1e"),
  2460 => (x"49",x"73",x"87",x"c6"),
  2461 => (x"71",x"29",x"b7",x"c8"),
  2462 => (x"fa",x"49",x"c1",x"1e"),
  2463 => (x"86",x"c8",x"87",x"fa"),
  2464 => (x"c2",x"87",x"c1",x"c6"),
  2465 => (x"4b",x"bf",x"ed",x"f8"),
  2466 => (x"87",x"dd",x"02",x"9b"),
  2467 => (x"bf",x"da",x"e1",x"c2"),
  2468 => (x"87",x"de",x"c7",x"49"),
  2469 => (x"c4",x"05",x"98",x"70"),
  2470 => (x"d2",x"4b",x"c0",x"87"),
  2471 => (x"49",x"e0",x"c2",x"87"),
  2472 => (x"c2",x"87",x"c3",x"c7"),
  2473 => (x"c6",x"58",x"de",x"e1"),
  2474 => (x"da",x"e1",x"c2",x"87"),
  2475 => (x"73",x"78",x"c0",x"48"),
  2476 => (x"05",x"99",x"c2",x"49"),
  2477 => (x"eb",x"c3",x"87",x"ce"),
  2478 => (x"d9",x"d6",x"ff",x"49"),
  2479 => (x"c2",x"49",x"70",x"87"),
  2480 => (x"87",x"c2",x"02",x"99"),
  2481 => (x"49",x"73",x"4c",x"fb"),
  2482 => (x"ce",x"05",x"99",x"c1"),
  2483 => (x"49",x"f4",x"c3",x"87"),
  2484 => (x"87",x"c2",x"d6",x"ff"),
  2485 => (x"99",x"c2",x"49",x"70"),
  2486 => (x"fa",x"87",x"c2",x"02"),
  2487 => (x"c8",x"49",x"73",x"4c"),
  2488 => (x"87",x"ce",x"05",x"99"),
  2489 => (x"ff",x"49",x"f5",x"c3"),
  2490 => (x"70",x"87",x"eb",x"d5"),
  2491 => (x"02",x"99",x"c2",x"49"),
  2492 => (x"f8",x"c2",x"87",x"d5"),
  2493 => (x"ca",x"02",x"bf",x"f5"),
  2494 => (x"88",x"c1",x"48",x"87"),
  2495 => (x"58",x"f9",x"f8",x"c2"),
  2496 => (x"ff",x"87",x"c2",x"c0"),
  2497 => (x"73",x"4d",x"c1",x"4c"),
  2498 => (x"05",x"99",x"c4",x"49"),
  2499 => (x"f2",x"c3",x"87",x"ce"),
  2500 => (x"c1",x"d5",x"ff",x"49"),
  2501 => (x"c2",x"49",x"70",x"87"),
  2502 => (x"87",x"dc",x"02",x"99"),
  2503 => (x"bf",x"f5",x"f8",x"c2"),
  2504 => (x"b7",x"c7",x"48",x"7e"),
  2505 => (x"cb",x"c0",x"03",x"a8"),
  2506 => (x"c1",x"48",x"6e",x"87"),
  2507 => (x"f9",x"f8",x"c2",x"80"),
  2508 => (x"87",x"c2",x"c0",x"58"),
  2509 => (x"4d",x"c1",x"4c",x"fe"),
  2510 => (x"ff",x"49",x"fd",x"c3"),
  2511 => (x"70",x"87",x"d7",x"d4"),
  2512 => (x"02",x"99",x"c2",x"49"),
  2513 => (x"c2",x"87",x"d5",x"c0"),
  2514 => (x"02",x"bf",x"f5",x"f8"),
  2515 => (x"c2",x"87",x"c9",x"c0"),
  2516 => (x"c0",x"48",x"f5",x"f8"),
  2517 => (x"87",x"c2",x"c0",x"78"),
  2518 => (x"4d",x"c1",x"4c",x"fd"),
  2519 => (x"ff",x"49",x"fa",x"c3"),
  2520 => (x"70",x"87",x"f3",x"d3"),
  2521 => (x"02",x"99",x"c2",x"49"),
  2522 => (x"c2",x"87",x"d9",x"c0"),
  2523 => (x"48",x"bf",x"f5",x"f8"),
  2524 => (x"03",x"a8",x"b7",x"c7"),
  2525 => (x"c2",x"87",x"c9",x"c0"),
  2526 => (x"c7",x"48",x"f5",x"f8"),
  2527 => (x"87",x"c2",x"c0",x"78"),
  2528 => (x"4d",x"c1",x"4c",x"fc"),
  2529 => (x"03",x"ac",x"b7",x"c0"),
  2530 => (x"c4",x"87",x"d1",x"c0"),
  2531 => (x"d8",x"c1",x"4a",x"66"),
  2532 => (x"c0",x"02",x"6a",x"82"),
  2533 => (x"4b",x"6a",x"87",x"c6"),
  2534 => (x"0f",x"73",x"49",x"74"),
  2535 => (x"f0",x"c3",x"1e",x"c0"),
  2536 => (x"49",x"da",x"c1",x"1e"),
  2537 => (x"c8",x"87",x"ce",x"f7"),
  2538 => (x"02",x"98",x"70",x"86"),
  2539 => (x"c8",x"87",x"e2",x"c0"),
  2540 => (x"f8",x"c2",x"48",x"a6"),
  2541 => (x"c8",x"78",x"bf",x"f5"),
  2542 => (x"91",x"cb",x"49",x"66"),
  2543 => (x"71",x"48",x"66",x"c4"),
  2544 => (x"6e",x"7e",x"70",x"80"),
  2545 => (x"c8",x"c0",x"02",x"bf"),
  2546 => (x"4b",x"bf",x"6e",x"87"),
  2547 => (x"73",x"49",x"66",x"c8"),
  2548 => (x"02",x"9d",x"75",x"0f"),
  2549 => (x"c2",x"87",x"c8",x"c0"),
  2550 => (x"49",x"bf",x"f5",x"f8"),
  2551 => (x"c2",x"87",x"fa",x"f2"),
  2552 => (x"02",x"bf",x"e2",x"e1"),
  2553 => (x"49",x"87",x"dd",x"c0"),
  2554 => (x"70",x"87",x"c7",x"c2"),
  2555 => (x"d3",x"c0",x"02",x"98"),
  2556 => (x"f5",x"f8",x"c2",x"87"),
  2557 => (x"e0",x"f2",x"49",x"bf"),
  2558 => (x"f4",x"49",x"c0",x"87"),
  2559 => (x"e1",x"c2",x"87",x"c0"),
  2560 => (x"78",x"c0",x"48",x"e2"),
  2561 => (x"da",x"f3",x"8e",x"f4"),
  2562 => (x"5b",x"5e",x"0e",x"87"),
  2563 => (x"1e",x"0e",x"5d",x"5c"),
  2564 => (x"f8",x"c2",x"4c",x"71"),
  2565 => (x"c1",x"49",x"bf",x"f1"),
  2566 => (x"c1",x"4d",x"a1",x"cd"),
  2567 => (x"7e",x"69",x"81",x"d1"),
  2568 => (x"cf",x"02",x"9c",x"74"),
  2569 => (x"4b",x"a5",x"c4",x"87"),
  2570 => (x"f8",x"c2",x"7b",x"74"),
  2571 => (x"f2",x"49",x"bf",x"f1"),
  2572 => (x"7b",x"6e",x"87",x"f9"),
  2573 => (x"c4",x"05",x"9c",x"74"),
  2574 => (x"c2",x"4b",x"c0",x"87"),
  2575 => (x"73",x"4b",x"c1",x"87"),
  2576 => (x"87",x"fa",x"f2",x"49"),
  2577 => (x"c7",x"02",x"66",x"d4"),
  2578 => (x"87",x"da",x"49",x"87"),
  2579 => (x"87",x"c2",x"4a",x"70"),
  2580 => (x"e1",x"c2",x"4a",x"c0"),
  2581 => (x"f2",x"26",x"5a",x"e6"),
  2582 => (x"00",x"00",x"87",x"c9"),
  2583 => (x"00",x"00",x"00",x"00"),
  2584 => (x"00",x"00",x"00",x"00"),
  2585 => (x"71",x"1e",x"00",x"00"),
  2586 => (x"bf",x"c8",x"ff",x"4a"),
  2587 => (x"48",x"a1",x"72",x"49"),
  2588 => (x"ff",x"1e",x"4f",x"26"),
  2589 => (x"fe",x"89",x"bf",x"c8"),
  2590 => (x"c0",x"c0",x"c0",x"c0"),
  2591 => (x"c4",x"01",x"a9",x"c0"),
  2592 => (x"c2",x"4a",x"c0",x"87"),
  2593 => (x"72",x"4a",x"c1",x"87"),
  2594 => (x"1e",x"4f",x"26",x"48"),
  2595 => (x"bf",x"d9",x"e3",x"c2"),
  2596 => (x"c2",x"b9",x"c1",x"49"),
  2597 => (x"ff",x"59",x"dd",x"e3"),
  2598 => (x"ff",x"c3",x"48",x"d4"),
  2599 => (x"48",x"d0",x"ff",x"78"),
  2600 => (x"ff",x"78",x"e1",x"c0"),
  2601 => (x"78",x"c1",x"48",x"d4"),
  2602 => (x"78",x"71",x"31",x"c4"),
  2603 => (x"c0",x"48",x"d0",x"ff"),
  2604 => (x"4f",x"26",x"78",x"e0"),
  2605 => (x"cd",x"e3",x"c2",x"1e"),
  2606 => (x"d8",x"f3",x"c2",x"1e"),
  2607 => (x"d1",x"fb",x"fd",x"49"),
  2608 => (x"70",x"86",x"c4",x"87"),
  2609 => (x"87",x"c3",x"02",x"98"),
  2610 => (x"26",x"87",x"c0",x"ff"),
  2611 => (x"4b",x"35",x"31",x"4f"),
  2612 => (x"20",x"20",x"5a",x"48"),
  2613 => (x"47",x"46",x"43",x"20"),
  2614 => (x"00",x"00",x"00",x"00"),
  2615 => (x"5b",x"5e",x"0e",x"00"),
  2616 => (x"c2",x"0e",x"5d",x"5c"),
  2617 => (x"4a",x"bf",x"e5",x"f8"),
  2618 => (x"bf",x"c6",x"e5",x"c2"),
  2619 => (x"bc",x"72",x"4c",x"49"),
  2620 => (x"c5",x"ff",x"4d",x"71"),
  2621 => (x"4b",x"c0",x"87",x"f7"),
  2622 => (x"99",x"d0",x"49",x"74"),
  2623 => (x"87",x"e7",x"c0",x"02"),
  2624 => (x"c8",x"48",x"d0",x"ff"),
  2625 => (x"d4",x"ff",x"78",x"e1"),
  2626 => (x"75",x"78",x"c5",x"48"),
  2627 => (x"02",x"99",x"d0",x"49"),
  2628 => (x"f0",x"c3",x"87",x"c3"),
  2629 => (x"f4",x"e5",x"c2",x"78"),
  2630 => (x"11",x"81",x"73",x"49"),
  2631 => (x"08",x"d4",x"ff",x"48"),
  2632 => (x"48",x"d0",x"ff",x"78"),
  2633 => (x"c1",x"78",x"e0",x"c0"),
  2634 => (x"c8",x"83",x"2d",x"2c"),
  2635 => (x"c7",x"ff",x"04",x"ab"),
  2636 => (x"f0",x"c4",x"ff",x"87"),
  2637 => (x"c6",x"e5",x"c2",x"87"),
  2638 => (x"e5",x"f8",x"c2",x"48"),
  2639 => (x"4d",x"26",x"78",x"bf"),
  2640 => (x"4b",x"26",x"4c",x"26"),
  2641 => (x"00",x"00",x"4f",x"26"),
  2642 => (x"c1",x"1e",x"00",x"00"),
  2643 => (x"de",x"48",x"d0",x"e7"),
  2644 => (x"dd",x"e5",x"c2",x"50"),
  2645 => (x"fa",x"d8",x"fe",x"49"),
  2646 => (x"26",x"48",x"c0",x"87"),
  2647 => (x"4f",x"54",x"4a",x"4f"),
  2648 => (x"55",x"52",x"54",x"55"),
  2649 => (x"43",x"52",x"41",x"4e"),
  2650 => (x"df",x"f2",x"1e",x"00"),
  2651 => (x"87",x"ed",x"fd",x"87"),
  2652 => (x"4f",x"26",x"87",x"f8"),
  2653 => (x"25",x"26",x"1e",x"16"),
  2654 => (x"3e",x"3d",x"36",x"2e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

