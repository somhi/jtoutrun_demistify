
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"44",x"4f",x"4d"),
     1 => (x"45",x"4d",x"41",x"4e"),
     2 => (x"46",x"45",x"44",x"00"),
     3 => (x"54",x"4c",x"55",x"41"),
     4 => (x"fa",x"00",x"30",x"3d"),
     5 => (x"00",x"00",x"00",x"1f"),
     6 => (x"04",x"00",x"00",x"20"),
     7 => (x"09",x"00",x"00",x"20"),
     8 => (x"1e",x"00",x"00",x"20"),
     9 => (x"c8",x"48",x"d0",x"ff"),
    10 => (x"48",x"71",x"78",x"c9"),
    11 => (x"78",x"08",x"d4",x"ff"),
    12 => (x"71",x"1e",x"4f",x"26"),
    13 => (x"87",x"eb",x"49",x"4a"),
    14 => (x"c8",x"48",x"d0",x"ff"),
    15 => (x"1e",x"4f",x"26",x"78"),
    16 => (x"4b",x"71",x"1e",x"73"),
    17 => (x"bf",x"fc",x"f9",x"c2"),
    18 => (x"c2",x"87",x"c3",x"02"),
    19 => (x"d0",x"ff",x"87",x"eb"),
    20 => (x"78",x"c9",x"c8",x"48"),
    21 => (x"e0",x"c0",x"49",x"73"),
    22 => (x"48",x"d4",x"ff",x"b1"),
    23 => (x"f9",x"c2",x"78",x"71"),
    24 => (x"78",x"c0",x"48",x"f0"),
    25 => (x"c5",x"02",x"66",x"c8"),
    26 => (x"49",x"ff",x"c3",x"87"),
    27 => (x"49",x"c0",x"87",x"c2"),
    28 => (x"59",x"f8",x"f9",x"c2"),
    29 => (x"c6",x"02",x"66",x"cc"),
    30 => (x"d5",x"d5",x"c5",x"87"),
    31 => (x"cf",x"87",x"c4",x"4a"),
    32 => (x"c2",x"4a",x"ff",x"ff"),
    33 => (x"c2",x"5a",x"fc",x"f9"),
    34 => (x"c1",x"48",x"fc",x"f9"),
    35 => (x"26",x"87",x"c4",x"78"),
    36 => (x"26",x"4c",x"26",x"4d"),
    37 => (x"0e",x"4f",x"26",x"4b"),
    38 => (x"5d",x"5c",x"5b",x"5e"),
    39 => (x"c2",x"4a",x"71",x"0e"),
    40 => (x"4c",x"bf",x"f8",x"f9"),
    41 => (x"cb",x"02",x"9a",x"72"),
    42 => (x"91",x"c8",x"49",x"87"),
    43 => (x"4b",x"f5",x"c0",x"c2"),
    44 => (x"87",x"c4",x"83",x"71"),
    45 => (x"4b",x"f5",x"c4",x"c2"),
    46 => (x"49",x"13",x"4d",x"c0"),
    47 => (x"f9",x"c2",x"99",x"74"),
    48 => (x"ff",x"b9",x"bf",x"f4"),
    49 => (x"78",x"71",x"48",x"d4"),
    50 => (x"85",x"2c",x"b7",x"c1"),
    51 => (x"04",x"ad",x"b7",x"c8"),
    52 => (x"f9",x"c2",x"87",x"e8"),
    53 => (x"c8",x"48",x"bf",x"f0"),
    54 => (x"f4",x"f9",x"c2",x"80"),
    55 => (x"87",x"ef",x"fe",x"58"),
    56 => (x"71",x"1e",x"73",x"1e"),
    57 => (x"9a",x"4a",x"13",x"4b"),
    58 => (x"72",x"87",x"cb",x"02"),
    59 => (x"87",x"e7",x"fe",x"49"),
    60 => (x"05",x"9a",x"4a",x"13"),
    61 => (x"da",x"fe",x"87",x"f5"),
    62 => (x"f9",x"c2",x"1e",x"87"),
    63 => (x"c2",x"49",x"bf",x"f0"),
    64 => (x"c1",x"48",x"f0",x"f9"),
    65 => (x"c0",x"c4",x"78",x"a1"),
    66 => (x"db",x"03",x"a9",x"b7"),
    67 => (x"48",x"d4",x"ff",x"87"),
    68 => (x"bf",x"f4",x"f9",x"c2"),
    69 => (x"f0",x"f9",x"c2",x"78"),
    70 => (x"f9",x"c2",x"49",x"bf"),
    71 => (x"a1",x"c1",x"48",x"f0"),
    72 => (x"b7",x"c0",x"c4",x"78"),
    73 => (x"87",x"e5",x"04",x"a9"),
    74 => (x"c8",x"48",x"d0",x"ff"),
    75 => (x"fc",x"f9",x"c2",x"78"),
    76 => (x"26",x"78",x"c0",x"48"),
    77 => (x"00",x"00",x"00",x"4f"),
    78 => (x"00",x"00",x"00",x"00"),
    79 => (x"00",x"00",x"00",x"00"),
    80 => (x"00",x"00",x"5f",x"5f"),
    81 => (x"03",x"03",x"00",x"00"),
    82 => (x"00",x"03",x"03",x"00"),
    83 => (x"7f",x"7f",x"14",x"00"),
    84 => (x"14",x"7f",x"7f",x"14"),
    85 => (x"2e",x"24",x"00",x"00"),
    86 => (x"12",x"3a",x"6b",x"6b"),
    87 => (x"36",x"6a",x"4c",x"00"),
    88 => (x"32",x"56",x"6c",x"18"),
    89 => (x"4f",x"7e",x"30",x"00"),
    90 => (x"68",x"3a",x"77",x"59"),
    91 => (x"04",x"00",x"00",x"40"),
    92 => (x"00",x"00",x"03",x"07"),
    93 => (x"1c",x"00",x"00",x"00"),
    94 => (x"00",x"41",x"63",x"3e"),
    95 => (x"41",x"00",x"00",x"00"),
    96 => (x"00",x"1c",x"3e",x"63"),
    97 => (x"3e",x"2a",x"08",x"00"),
    98 => (x"2a",x"3e",x"1c",x"1c"),
    99 => (x"08",x"08",x"00",x"08"),
   100 => (x"08",x"08",x"3e",x"3e"),
   101 => (x"80",x"00",x"00",x"00"),
   102 => (x"00",x"00",x"60",x"e0"),
   103 => (x"08",x"08",x"00",x"00"),
   104 => (x"08",x"08",x"08",x"08"),
   105 => (x"00",x"00",x"00",x"00"),
   106 => (x"00",x"00",x"60",x"60"),
   107 => (x"30",x"60",x"40",x"00"),
   108 => (x"03",x"06",x"0c",x"18"),
   109 => (x"7f",x"3e",x"00",x"01"),
   110 => (x"3e",x"7f",x"4d",x"59"),
   111 => (x"06",x"04",x"00",x"00"),
   112 => (x"00",x"00",x"7f",x"7f"),
   113 => (x"63",x"42",x"00",x"00"),
   114 => (x"46",x"4f",x"59",x"71"),
   115 => (x"63",x"22",x"00",x"00"),
   116 => (x"36",x"7f",x"49",x"49"),
   117 => (x"16",x"1c",x"18",x"00"),
   118 => (x"10",x"7f",x"7f",x"13"),
   119 => (x"67",x"27",x"00",x"00"),
   120 => (x"39",x"7d",x"45",x"45"),
   121 => (x"7e",x"3c",x"00",x"00"),
   122 => (x"30",x"79",x"49",x"4b"),
   123 => (x"01",x"01",x"00",x"00"),
   124 => (x"07",x"0f",x"79",x"71"),
   125 => (x"7f",x"36",x"00",x"00"),
   126 => (x"36",x"7f",x"49",x"49"),
   127 => (x"4f",x"06",x"00",x"00"),
   128 => (x"1e",x"3f",x"69",x"49"),
   129 => (x"00",x"00",x"00",x"00"),
   130 => (x"00",x"00",x"66",x"66"),
   131 => (x"80",x"00",x"00",x"00"),
   132 => (x"00",x"00",x"66",x"e6"),
   133 => (x"08",x"08",x"00",x"00"),
   134 => (x"22",x"22",x"14",x"14"),
   135 => (x"14",x"14",x"00",x"00"),
   136 => (x"14",x"14",x"14",x"14"),
   137 => (x"22",x"22",x"00",x"00"),
   138 => (x"08",x"08",x"14",x"14"),
   139 => (x"03",x"02",x"00",x"00"),
   140 => (x"06",x"0f",x"59",x"51"),
   141 => (x"41",x"7f",x"3e",x"00"),
   142 => (x"1e",x"1f",x"55",x"5d"),
   143 => (x"7f",x"7e",x"00",x"00"),
   144 => (x"7e",x"7f",x"09",x"09"),
   145 => (x"7f",x"7f",x"00",x"00"),
   146 => (x"36",x"7f",x"49",x"49"),
   147 => (x"3e",x"1c",x"00",x"00"),
   148 => (x"41",x"41",x"41",x"63"),
   149 => (x"7f",x"7f",x"00",x"00"),
   150 => (x"1c",x"3e",x"63",x"41"),
   151 => (x"7f",x"7f",x"00",x"00"),
   152 => (x"41",x"41",x"49",x"49"),
   153 => (x"7f",x"7f",x"00",x"00"),
   154 => (x"01",x"01",x"09",x"09"),
   155 => (x"7f",x"3e",x"00",x"00"),
   156 => (x"7a",x"7b",x"49",x"41"),
   157 => (x"7f",x"7f",x"00",x"00"),
   158 => (x"7f",x"7f",x"08",x"08"),
   159 => (x"41",x"00",x"00",x"00"),
   160 => (x"00",x"41",x"7f",x"7f"),
   161 => (x"60",x"20",x"00",x"00"),
   162 => (x"3f",x"7f",x"40",x"40"),
   163 => (x"08",x"7f",x"7f",x"00"),
   164 => (x"41",x"63",x"36",x"1c"),
   165 => (x"7f",x"7f",x"00",x"00"),
   166 => (x"40",x"40",x"40",x"40"),
   167 => (x"06",x"7f",x"7f",x"00"),
   168 => (x"7f",x"7f",x"06",x"0c"),
   169 => (x"06",x"7f",x"7f",x"00"),
   170 => (x"7f",x"7f",x"18",x"0c"),
   171 => (x"7f",x"3e",x"00",x"00"),
   172 => (x"3e",x"7f",x"41",x"41"),
   173 => (x"7f",x"7f",x"00",x"00"),
   174 => (x"06",x"0f",x"09",x"09"),
   175 => (x"41",x"7f",x"3e",x"00"),
   176 => (x"40",x"7e",x"7f",x"61"),
   177 => (x"7f",x"7f",x"00",x"00"),
   178 => (x"66",x"7f",x"19",x"09"),
   179 => (x"6f",x"26",x"00",x"00"),
   180 => (x"32",x"7b",x"59",x"4d"),
   181 => (x"01",x"01",x"00",x"00"),
   182 => (x"01",x"01",x"7f",x"7f"),
   183 => (x"7f",x"3f",x"00",x"00"),
   184 => (x"3f",x"7f",x"40",x"40"),
   185 => (x"3f",x"0f",x"00",x"00"),
   186 => (x"0f",x"3f",x"70",x"70"),
   187 => (x"30",x"7f",x"7f",x"00"),
   188 => (x"7f",x"7f",x"30",x"18"),
   189 => (x"36",x"63",x"41",x"00"),
   190 => (x"63",x"36",x"1c",x"1c"),
   191 => (x"06",x"03",x"01",x"41"),
   192 => (x"03",x"06",x"7c",x"7c"),
   193 => (x"59",x"71",x"61",x"01"),
   194 => (x"41",x"43",x"47",x"4d"),
   195 => (x"7f",x"00",x"00",x"00"),
   196 => (x"00",x"41",x"41",x"7f"),
   197 => (x"06",x"03",x"01",x"00"),
   198 => (x"60",x"30",x"18",x"0c"),
   199 => (x"41",x"00",x"00",x"40"),
   200 => (x"00",x"7f",x"7f",x"41"),
   201 => (x"06",x"0c",x"08",x"00"),
   202 => (x"08",x"0c",x"06",x"03"),
   203 => (x"80",x"80",x"80",x"00"),
   204 => (x"80",x"80",x"80",x"80"),
   205 => (x"00",x"00",x"00",x"00"),
   206 => (x"00",x"04",x"07",x"03"),
   207 => (x"74",x"20",x"00",x"00"),
   208 => (x"78",x"7c",x"54",x"54"),
   209 => (x"7f",x"7f",x"00",x"00"),
   210 => (x"38",x"7c",x"44",x"44"),
   211 => (x"7c",x"38",x"00",x"00"),
   212 => (x"00",x"44",x"44",x"44"),
   213 => (x"7c",x"38",x"00",x"00"),
   214 => (x"7f",x"7f",x"44",x"44"),
   215 => (x"7c",x"38",x"00",x"00"),
   216 => (x"18",x"5c",x"54",x"54"),
   217 => (x"7e",x"04",x"00",x"00"),
   218 => (x"00",x"05",x"05",x"7f"),
   219 => (x"bc",x"18",x"00",x"00"),
   220 => (x"7c",x"fc",x"a4",x"a4"),
   221 => (x"7f",x"7f",x"00",x"00"),
   222 => (x"78",x"7c",x"04",x"04"),
   223 => (x"00",x"00",x"00",x"00"),
   224 => (x"00",x"40",x"7d",x"3d"),
   225 => (x"80",x"80",x"00",x"00"),
   226 => (x"00",x"7d",x"fd",x"80"),
   227 => (x"7f",x"7f",x"00",x"00"),
   228 => (x"44",x"6c",x"38",x"10"),
   229 => (x"00",x"00",x"00",x"00"),
   230 => (x"00",x"40",x"7f",x"3f"),
   231 => (x"0c",x"7c",x"7c",x"00"),
   232 => (x"78",x"7c",x"0c",x"18"),
   233 => (x"7c",x"7c",x"00",x"00"),
   234 => (x"78",x"7c",x"04",x"04"),
   235 => (x"7c",x"38",x"00",x"00"),
   236 => (x"38",x"7c",x"44",x"44"),
   237 => (x"fc",x"fc",x"00",x"00"),
   238 => (x"18",x"3c",x"24",x"24"),
   239 => (x"3c",x"18",x"00",x"00"),
   240 => (x"fc",x"fc",x"24",x"24"),
   241 => (x"7c",x"7c",x"00",x"00"),
   242 => (x"08",x"0c",x"04",x"04"),
   243 => (x"5c",x"48",x"00",x"00"),
   244 => (x"20",x"74",x"54",x"54"),
   245 => (x"3f",x"04",x"00",x"00"),
   246 => (x"00",x"44",x"44",x"7f"),
   247 => (x"7c",x"3c",x"00",x"00"),
   248 => (x"7c",x"7c",x"40",x"40"),
   249 => (x"3c",x"1c",x"00",x"00"),
   250 => (x"1c",x"3c",x"60",x"60"),
   251 => (x"60",x"7c",x"3c",x"00"),
   252 => (x"3c",x"7c",x"60",x"30"),
   253 => (x"38",x"6c",x"44",x"00"),
   254 => (x"44",x"6c",x"38",x"10"),
   255 => (x"bc",x"1c",x"00",x"00"),
   256 => (x"1c",x"3c",x"60",x"e0"),
   257 => (x"64",x"44",x"00",x"00"),
   258 => (x"44",x"4c",x"5c",x"74"),
   259 => (x"08",x"08",x"00",x"00"),
   260 => (x"41",x"41",x"77",x"3e"),
   261 => (x"00",x"00",x"00",x"00"),
   262 => (x"00",x"00",x"7f",x"7f"),
   263 => (x"41",x"41",x"00",x"00"),
   264 => (x"08",x"08",x"3e",x"77"),
   265 => (x"01",x"01",x"02",x"00"),
   266 => (x"01",x"02",x"02",x"03"),
   267 => (x"7f",x"7f",x"7f",x"00"),
   268 => (x"7f",x"7f",x"7f",x"7f"),
   269 => (x"1c",x"08",x"08",x"00"),
   270 => (x"7f",x"3e",x"3e",x"1c"),
   271 => (x"3e",x"7f",x"7f",x"7f"),
   272 => (x"08",x"1c",x"1c",x"3e"),
   273 => (x"18",x"10",x"00",x"08"),
   274 => (x"10",x"18",x"7c",x"7c"),
   275 => (x"30",x"10",x"00",x"00"),
   276 => (x"10",x"30",x"7c",x"7c"),
   277 => (x"60",x"30",x"10",x"00"),
   278 => (x"06",x"1e",x"78",x"60"),
   279 => (x"3c",x"66",x"42",x"00"),
   280 => (x"42",x"66",x"3c",x"18"),
   281 => (x"6a",x"38",x"78",x"00"),
   282 => (x"38",x"6c",x"c6",x"c2"),
   283 => (x"00",x"00",x"60",x"00"),
   284 => (x"60",x"00",x"00",x"60"),
   285 => (x"5b",x"5e",x"0e",x"00"),
   286 => (x"1e",x"0e",x"5d",x"5c"),
   287 => (x"fa",x"c2",x"4c",x"71"),
   288 => (x"c0",x"4d",x"bf",x"cd"),
   289 => (x"74",x"1e",x"c0",x"4b"),
   290 => (x"87",x"c7",x"02",x"ab"),
   291 => (x"c0",x"48",x"a6",x"c4"),
   292 => (x"c4",x"87",x"c5",x"78"),
   293 => (x"78",x"c1",x"48",x"a6"),
   294 => (x"73",x"1e",x"66",x"c4"),
   295 => (x"87",x"df",x"ee",x"49"),
   296 => (x"e0",x"c0",x"86",x"c8"),
   297 => (x"87",x"ef",x"ef",x"49"),
   298 => (x"6a",x"4a",x"a5",x"c4"),
   299 => (x"87",x"f0",x"f0",x"49"),
   300 => (x"cb",x"87",x"c6",x"f1"),
   301 => (x"c8",x"83",x"c1",x"85"),
   302 => (x"ff",x"04",x"ab",x"b7"),
   303 => (x"26",x"26",x"87",x"c7"),
   304 => (x"26",x"4c",x"26",x"4d"),
   305 => (x"1e",x"4f",x"26",x"4b"),
   306 => (x"fa",x"c2",x"4a",x"71"),
   307 => (x"fa",x"c2",x"5a",x"d1"),
   308 => (x"78",x"c7",x"48",x"d1"),
   309 => (x"87",x"dd",x"fe",x"49"),
   310 => (x"73",x"1e",x"4f",x"26"),
   311 => (x"c0",x"4a",x"71",x"1e"),
   312 => (x"d3",x"03",x"aa",x"b7"),
   313 => (x"fa",x"e0",x"c2",x"87"),
   314 => (x"87",x"c4",x"05",x"bf"),
   315 => (x"87",x"c2",x"4b",x"c1"),
   316 => (x"e0",x"c2",x"4b",x"c0"),
   317 => (x"87",x"c4",x"5b",x"fe"),
   318 => (x"5a",x"fe",x"e0",x"c2"),
   319 => (x"bf",x"fa",x"e0",x"c2"),
   320 => (x"c1",x"9a",x"c1",x"4a"),
   321 => (x"ec",x"49",x"a2",x"c0"),
   322 => (x"48",x"fc",x"87",x"e8"),
   323 => (x"bf",x"fa",x"e0",x"c2"),
   324 => (x"87",x"ef",x"fe",x"78"),
   325 => (x"c4",x"4a",x"71",x"1e"),
   326 => (x"49",x"72",x"1e",x"66"),
   327 => (x"87",x"dd",x"df",x"ff"),
   328 => (x"1e",x"4f",x"26",x"26"),
   329 => (x"bf",x"fa",x"e0",x"c2"),
   330 => (x"cd",x"dc",x"ff",x"49"),
   331 => (x"c5",x"fa",x"c2",x"87"),
   332 => (x"78",x"bf",x"e8",x"48"),
   333 => (x"48",x"c1",x"fa",x"c2"),
   334 => (x"c2",x"78",x"bf",x"ec"),
   335 => (x"4a",x"bf",x"c5",x"fa"),
   336 => (x"99",x"ff",x"c3",x"49"),
   337 => (x"72",x"2a",x"b7",x"c8"),
   338 => (x"c2",x"b0",x"71",x"48"),
   339 => (x"26",x"58",x"cd",x"fa"),
   340 => (x"5b",x"5e",x"0e",x"4f"),
   341 => (x"71",x"0e",x"5d",x"5c"),
   342 => (x"87",x"c7",x"ff",x"4b"),
   343 => (x"48",x"c0",x"fa",x"c2"),
   344 => (x"49",x"73",x"50",x"c0"),
   345 => (x"87",x"f2",x"db",x"ff"),
   346 => (x"c2",x"4c",x"49",x"70"),
   347 => (x"49",x"ee",x"cb",x"9c"),
   348 => (x"70",x"87",x"cf",x"cb"),
   349 => (x"fa",x"c2",x"4d",x"49"),
   350 => (x"05",x"bf",x"97",x"c0"),
   351 => (x"d0",x"87",x"e4",x"c1"),
   352 => (x"fa",x"c2",x"49",x"66"),
   353 => (x"05",x"99",x"bf",x"c9"),
   354 => (x"66",x"d4",x"87",x"d7"),
   355 => (x"c1",x"fa",x"c2",x"49"),
   356 => (x"cc",x"05",x"99",x"bf"),
   357 => (x"ff",x"49",x"73",x"87"),
   358 => (x"70",x"87",x"ff",x"da"),
   359 => (x"c2",x"c1",x"02",x"98"),
   360 => (x"fd",x"4c",x"c1",x"87"),
   361 => (x"49",x"75",x"87",x"fd"),
   362 => (x"70",x"87",x"e3",x"ca"),
   363 => (x"87",x"c6",x"02",x"98"),
   364 => (x"48",x"c0",x"fa",x"c2"),
   365 => (x"fa",x"c2",x"50",x"c1"),
   366 => (x"05",x"bf",x"97",x"c0"),
   367 => (x"c2",x"87",x"e4",x"c0"),
   368 => (x"49",x"bf",x"c9",x"fa"),
   369 => (x"05",x"99",x"66",x"d0"),
   370 => (x"c2",x"87",x"d6",x"ff"),
   371 => (x"49",x"bf",x"c1",x"fa"),
   372 => (x"05",x"99",x"66",x"d4"),
   373 => (x"73",x"87",x"ca",x"ff"),
   374 => (x"fd",x"d9",x"ff",x"49"),
   375 => (x"05",x"98",x"70",x"87"),
   376 => (x"74",x"87",x"fe",x"fe"),
   377 => (x"87",x"d7",x"fb",x"48"),
   378 => (x"5c",x"5b",x"5e",x"0e"),
   379 => (x"86",x"f4",x"0e",x"5d"),
   380 => (x"ec",x"4c",x"4d",x"c0"),
   381 => (x"a6",x"c4",x"7e",x"bf"),
   382 => (x"cd",x"fa",x"c2",x"48"),
   383 => (x"1e",x"c1",x"78",x"bf"),
   384 => (x"49",x"c7",x"1e",x"c0"),
   385 => (x"c8",x"87",x"ca",x"fd"),
   386 => (x"02",x"98",x"70",x"86"),
   387 => (x"49",x"ff",x"87",x"ce"),
   388 => (x"c1",x"87",x"c7",x"fb"),
   389 => (x"d9",x"ff",x"49",x"da"),
   390 => (x"4d",x"c1",x"87",x"c0"),
   391 => (x"97",x"c0",x"fa",x"c2"),
   392 => (x"87",x"c3",x"02",x"bf"),
   393 => (x"c2",x"87",x"c0",x"c9"),
   394 => (x"4b",x"bf",x"c5",x"fa"),
   395 => (x"bf",x"fa",x"e0",x"c2"),
   396 => (x"87",x"eb",x"c0",x"05"),
   397 => (x"ff",x"49",x"fd",x"c3"),
   398 => (x"c3",x"87",x"df",x"d8"),
   399 => (x"d8",x"ff",x"49",x"fa"),
   400 => (x"49",x"73",x"87",x"d8"),
   401 => (x"71",x"99",x"ff",x"c3"),
   402 => (x"fb",x"49",x"c0",x"1e"),
   403 => (x"49",x"73",x"87",x"c6"),
   404 => (x"71",x"29",x"b7",x"c8"),
   405 => (x"fa",x"49",x"c1",x"1e"),
   406 => (x"86",x"c8",x"87",x"fa"),
   407 => (x"c2",x"87",x"c1",x"c6"),
   408 => (x"4b",x"bf",x"c9",x"fa"),
   409 => (x"87",x"dd",x"02",x"9b"),
   410 => (x"bf",x"f6",x"e0",x"c2"),
   411 => (x"87",x"de",x"c7",x"49"),
   412 => (x"c4",x"05",x"98",x"70"),
   413 => (x"d2",x"4b",x"c0",x"87"),
   414 => (x"49",x"e0",x"c2",x"87"),
   415 => (x"c2",x"87",x"c3",x"c7"),
   416 => (x"c6",x"58",x"fa",x"e0"),
   417 => (x"f6",x"e0",x"c2",x"87"),
   418 => (x"73",x"78",x"c0",x"48"),
   419 => (x"05",x"99",x"c2",x"49"),
   420 => (x"eb",x"c3",x"87",x"ce"),
   421 => (x"c1",x"d7",x"ff",x"49"),
   422 => (x"c2",x"49",x"70",x"87"),
   423 => (x"87",x"c2",x"02",x"99"),
   424 => (x"49",x"73",x"4c",x"fb"),
   425 => (x"ce",x"05",x"99",x"c1"),
   426 => (x"49",x"f4",x"c3",x"87"),
   427 => (x"87",x"ea",x"d6",x"ff"),
   428 => (x"99",x"c2",x"49",x"70"),
   429 => (x"fa",x"87",x"c2",x"02"),
   430 => (x"c8",x"49",x"73",x"4c"),
   431 => (x"87",x"ce",x"05",x"99"),
   432 => (x"ff",x"49",x"f5",x"c3"),
   433 => (x"70",x"87",x"d3",x"d6"),
   434 => (x"02",x"99",x"c2",x"49"),
   435 => (x"fa",x"c2",x"87",x"d5"),
   436 => (x"ca",x"02",x"bf",x"d1"),
   437 => (x"88",x"c1",x"48",x"87"),
   438 => (x"58",x"d5",x"fa",x"c2"),
   439 => (x"ff",x"87",x"c2",x"c0"),
   440 => (x"73",x"4d",x"c1",x"4c"),
   441 => (x"05",x"99",x"c4",x"49"),
   442 => (x"f2",x"c3",x"87",x"ce"),
   443 => (x"e9",x"d5",x"ff",x"49"),
   444 => (x"c2",x"49",x"70",x"87"),
   445 => (x"87",x"dc",x"02",x"99"),
   446 => (x"bf",x"d1",x"fa",x"c2"),
   447 => (x"b7",x"c7",x"48",x"7e"),
   448 => (x"cb",x"c0",x"03",x"a8"),
   449 => (x"c1",x"48",x"6e",x"87"),
   450 => (x"d5",x"fa",x"c2",x"80"),
   451 => (x"87",x"c2",x"c0",x"58"),
   452 => (x"4d",x"c1",x"4c",x"fe"),
   453 => (x"ff",x"49",x"fd",x"c3"),
   454 => (x"70",x"87",x"ff",x"d4"),
   455 => (x"02",x"99",x"c2",x"49"),
   456 => (x"c2",x"87",x"d5",x"c0"),
   457 => (x"02",x"bf",x"d1",x"fa"),
   458 => (x"c2",x"87",x"c9",x"c0"),
   459 => (x"c0",x"48",x"d1",x"fa"),
   460 => (x"87",x"c2",x"c0",x"78"),
   461 => (x"4d",x"c1",x"4c",x"fd"),
   462 => (x"ff",x"49",x"fa",x"c3"),
   463 => (x"70",x"87",x"db",x"d4"),
   464 => (x"02",x"99",x"c2",x"49"),
   465 => (x"c2",x"87",x"d9",x"c0"),
   466 => (x"48",x"bf",x"d1",x"fa"),
   467 => (x"03",x"a8",x"b7",x"c7"),
   468 => (x"c2",x"87",x"c9",x"c0"),
   469 => (x"c7",x"48",x"d1",x"fa"),
   470 => (x"87",x"c2",x"c0",x"78"),
   471 => (x"4d",x"c1",x"4c",x"fc"),
   472 => (x"03",x"ac",x"b7",x"c0"),
   473 => (x"c4",x"87",x"d1",x"c0"),
   474 => (x"d8",x"c1",x"4a",x"66"),
   475 => (x"c0",x"02",x"6a",x"82"),
   476 => (x"4b",x"6a",x"87",x"c6"),
   477 => (x"0f",x"73",x"49",x"74"),
   478 => (x"f0",x"c3",x"1e",x"c0"),
   479 => (x"49",x"da",x"c1",x"1e"),
   480 => (x"c8",x"87",x"ce",x"f7"),
   481 => (x"02",x"98",x"70",x"86"),
   482 => (x"c8",x"87",x"e2",x"c0"),
   483 => (x"fa",x"c2",x"48",x"a6"),
   484 => (x"c8",x"78",x"bf",x"d1"),
   485 => (x"91",x"cb",x"49",x"66"),
   486 => (x"71",x"48",x"66",x"c4"),
   487 => (x"6e",x"7e",x"70",x"80"),
   488 => (x"c8",x"c0",x"02",x"bf"),
   489 => (x"4b",x"bf",x"6e",x"87"),
   490 => (x"73",x"49",x"66",x"c8"),
   491 => (x"02",x"9d",x"75",x"0f"),
   492 => (x"c2",x"87",x"c8",x"c0"),
   493 => (x"49",x"bf",x"d1",x"fa"),
   494 => (x"c2",x"87",x"fa",x"f2"),
   495 => (x"02",x"bf",x"fe",x"e0"),
   496 => (x"49",x"87",x"dd",x"c0"),
   497 => (x"70",x"87",x"c7",x"c2"),
   498 => (x"d3",x"c0",x"02",x"98"),
   499 => (x"d1",x"fa",x"c2",x"87"),
   500 => (x"e0",x"f2",x"49",x"bf"),
   501 => (x"f4",x"49",x"c0",x"87"),
   502 => (x"e0",x"c2",x"87",x"c0"),
   503 => (x"78",x"c0",x"48",x"fe"),
   504 => (x"da",x"f3",x"8e",x"f4"),
   505 => (x"5b",x"5e",x"0e",x"87"),
   506 => (x"1e",x"0e",x"5d",x"5c"),
   507 => (x"fa",x"c2",x"4c",x"71"),
   508 => (x"c1",x"49",x"bf",x"cd"),
   509 => (x"c1",x"4d",x"a1",x"cd"),
   510 => (x"7e",x"69",x"81",x"d1"),
   511 => (x"cf",x"02",x"9c",x"74"),
   512 => (x"4b",x"a5",x"c4",x"87"),
   513 => (x"fa",x"c2",x"7b",x"74"),
   514 => (x"f2",x"49",x"bf",x"cd"),
   515 => (x"7b",x"6e",x"87",x"f9"),
   516 => (x"c4",x"05",x"9c",x"74"),
   517 => (x"c2",x"4b",x"c0",x"87"),
   518 => (x"73",x"4b",x"c1",x"87"),
   519 => (x"87",x"fa",x"f2",x"49"),
   520 => (x"c7",x"02",x"66",x"d4"),
   521 => (x"87",x"da",x"49",x"87"),
   522 => (x"87",x"c2",x"4a",x"70"),
   523 => (x"e1",x"c2",x"4a",x"c0"),
   524 => (x"f2",x"26",x"5a",x"c2"),
   525 => (x"00",x"00",x"87",x"c9"),
   526 => (x"00",x"00",x"00",x"00"),
   527 => (x"00",x"00",x"00",x"00"),
   528 => (x"71",x"1e",x"00",x"00"),
   529 => (x"bf",x"c8",x"ff",x"4a"),
   530 => (x"48",x"a1",x"72",x"49"),
   531 => (x"ff",x"1e",x"4f",x"26"),
   532 => (x"fe",x"89",x"bf",x"c8"),
   533 => (x"c0",x"c0",x"c0",x"c0"),
   534 => (x"c4",x"01",x"a9",x"c0"),
   535 => (x"c2",x"4a",x"c0",x"87"),
   536 => (x"72",x"4a",x"c1",x"87"),
   537 => (x"1e",x"4f",x"26",x"48"),
   538 => (x"bf",x"f5",x"e2",x"c2"),
   539 => (x"c2",x"b9",x"c1",x"49"),
   540 => (x"ff",x"59",x"f9",x"e2"),
   541 => (x"ff",x"c3",x"48",x"d4"),
   542 => (x"48",x"d0",x"ff",x"78"),
   543 => (x"ff",x"78",x"e1",x"c0"),
   544 => (x"78",x"c1",x"48",x"d4"),
   545 => (x"78",x"71",x"31",x"c4"),
   546 => (x"c0",x"48",x"d0",x"ff"),
   547 => (x"4f",x"26",x"78",x"e0"),
   548 => (x"e9",x"e2",x"c2",x"1e"),
   549 => (x"f4",x"f4",x"c2",x"1e"),
   550 => (x"d4",x"fd",x"fd",x"49"),
   551 => (x"70",x"86",x"c4",x"87"),
   552 => (x"87",x"c3",x"02",x"98"),
   553 => (x"26",x"87",x"c0",x"ff"),
   554 => (x"4b",x"35",x"31",x"4f"),
   555 => (x"20",x"20",x"5a",x"48"),
   556 => (x"47",x"46",x"43",x"20"),
   557 => (x"00",x"00",x"00",x"00"),
   558 => (x"5b",x"5e",x"0e",x"00"),
   559 => (x"c2",x"0e",x"5d",x"5c"),
   560 => (x"4a",x"bf",x"c1",x"fa"),
   561 => (x"bf",x"e2",x"e4",x"c2"),
   562 => (x"bc",x"72",x"4c",x"49"),
   563 => (x"c6",x"ff",x"4d",x"71"),
   564 => (x"4b",x"c0",x"87",x"de"),
   565 => (x"99",x"d0",x"49",x"74"),
   566 => (x"87",x"e7",x"c0",x"02"),
   567 => (x"c8",x"48",x"d0",x"ff"),
   568 => (x"d4",x"ff",x"78",x"e1"),
   569 => (x"75",x"78",x"c5",x"48"),
   570 => (x"02",x"99",x"d0",x"49"),
   571 => (x"f0",x"c3",x"87",x"c3"),
   572 => (x"cf",x"e7",x"c2",x"78"),
   573 => (x"11",x"81",x"73",x"49"),
   574 => (x"08",x"d4",x"ff",x"48"),
   575 => (x"48",x"d0",x"ff",x"78"),
   576 => (x"c1",x"78",x"e0",x"c0"),
   577 => (x"c8",x"83",x"2d",x"2c"),
   578 => (x"c7",x"ff",x"04",x"ab"),
   579 => (x"d7",x"c5",x"ff",x"87"),
   580 => (x"e2",x"e4",x"c2",x"87"),
   581 => (x"c1",x"fa",x"c2",x"48"),
   582 => (x"4d",x"26",x"78",x"bf"),
   583 => (x"4b",x"26",x"4c",x"26"),
   584 => (x"00",x"00",x"4f",x"26"),
   585 => (x"73",x"1e",x"00",x"00"),
   586 => (x"c1",x"4b",x"c0",x"1e"),
   587 => (x"de",x"48",x"d7",x"e7"),
   588 => (x"c2",x"1e",x"c8",x"50"),
   589 => (x"fe",x"49",x"d5",x"fa"),
   590 => (x"c4",x"87",x"c1",x"d5"),
   591 => (x"c2",x"1e",x"72",x"86"),
   592 => (x"c2",x"48",x"d8",x"e6"),
   593 => (x"c4",x"49",x"dd",x"fa"),
   594 => (x"41",x"20",x"4a",x"a1"),
   595 => (x"f9",x"05",x"aa",x"71"),
   596 => (x"c2",x"4a",x"26",x"87"),
   597 => (x"fd",x"49",x"dc",x"e6"),
   598 => (x"70",x"87",x"f7",x"f8"),
   599 => (x"c5",x"02",x"9a",x"4a"),
   600 => (x"c7",x"fe",x"49",x"87"),
   601 => (x"1e",x"72",x"87",x"e0"),
   602 => (x"48",x"e8",x"e6",x"c2"),
   603 => (x"49",x"dd",x"fa",x"c2"),
   604 => (x"20",x"4a",x"a1",x"c4"),
   605 => (x"05",x"aa",x"71",x"41"),
   606 => (x"4a",x"26",x"87",x"f9"),
   607 => (x"49",x"d5",x"fa",x"c2"),
   608 => (x"87",x"d1",x"d9",x"fe"),
   609 => (x"c4",x"05",x"98",x"70"),
   610 => (x"ec",x"e6",x"c2",x"87"),
   611 => (x"fe",x"49",x"c0",x"4b"),
   612 => (x"73",x"87",x"d5",x"c5"),
   613 => (x"87",x"c6",x"fe",x"48"),
   614 => (x"00",x"20",x"20",x"20"),
   615 => (x"45",x"54",x"4f",x"4a"),
   616 => (x"20",x"20",x"4f",x"47"),
   617 => (x"00",x"20",x"20",x"20"),
   618 => (x"00",x"43",x"52",x"41"),
   619 => (x"20",x"43",x"52",x"41"),
   620 => (x"20",x"74",x"6f",x"6e"),
   621 => (x"6e",x"75",x"6f",x"66"),
   622 => (x"4c",x"20",x"2e",x"64"),
   623 => (x"20",x"64",x"61",x"6f"),
   624 => (x"00",x"43",x"52",x"41"),
   625 => (x"87",x"e0",x"f0",x"1e"),
   626 => (x"f8",x"87",x"ee",x"fb"),
   627 => (x"16",x"4f",x"26",x"87"),
   628 => (x"2e",x"25",x"26",x"1e"),
   629 => (x"2e",x"3e",x"3d",x"36"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

