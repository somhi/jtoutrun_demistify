library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fcf7c287",
    12 => x"86c0c84e",
    13 => x"49fcf7c2",
    14 => x"48fce4c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e6e5",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"8148731e",
    47 => x"7205a973",
    48 => x"2687f953",
    49 => x"4a711e4f",
    50 => x"484966c4",
    51 => x"a6c888c1",
    52 => x"02997158",
    53 => x"d4ff87d6",
    54 => x"78ffc348",
    55 => x"66c45268",
    56 => x"88c14849",
    57 => x"7158a6c8",
    58 => x"87ea0599",
    59 => x"731e4f26",
    60 => x"4bd4ff1e",
    61 => x"6b7bffc3",
    62 => x"7bffc34a",
    63 => x"32c8496b",
    64 => x"ffc3b172",
    65 => x"c84a6b7b",
    66 => x"c3b27131",
    67 => x"496b7bff",
    68 => x"b17232c8",
    69 => x"87c44871",
    70 => x"4c264d26",
    71 => x"4f264b26",
    72 => x"5c5b5e0e",
    73 => x"4a710e5d",
    74 => x"724cd4ff",
    75 => x"99ffc349",
    76 => x"e4c27c71",
    77 => x"c805bffc",
    78 => x"4866d087",
    79 => x"a6d430c9",
    80 => x"4966d058",
    81 => x"ffc329d8",
    82 => x"d07c7199",
    83 => x"29d04966",
    84 => x"7199ffc3",
    85 => x"4966d07c",
    86 => x"ffc329c8",
    87 => x"d07c7199",
    88 => x"ffc34966",
    89 => x"727c7199",
    90 => x"c329d049",
    91 => x"7c7199ff",
    92 => x"f0c94b6c",
    93 => x"ffc34dff",
    94 => x"87d005ab",
    95 => x"6c7cffc3",
    96 => x"028dc14b",
    97 => x"ffc387c6",
    98 => x"87f002ab",
    99 => x"c7fe4873",
   100 => x"49c01e87",
   101 => x"c348d4ff",
   102 => x"81c178ff",
   103 => x"a9b7c8c3",
   104 => x"2687f104",
   105 => x"1e731e4f",
   106 => x"f8c487e7",
   107 => x"1ec04bdf",
   108 => x"c1f0ffc0",
   109 => x"e7fd49f7",
   110 => x"c186c487",
   111 => x"eac005a8",
   112 => x"48d4ff87",
   113 => x"c178ffc3",
   114 => x"c0c0c0c0",
   115 => x"e1c01ec0",
   116 => x"49e9c1f0",
   117 => x"c487c9fd",
   118 => x"05987086",
   119 => x"d4ff87ca",
   120 => x"78ffc348",
   121 => x"87cb48c1",
   122 => x"c187e6fe",
   123 => x"fdfe058b",
   124 => x"fc48c087",
   125 => x"731e87e6",
   126 => x"48d4ff1e",
   127 => x"d378ffc3",
   128 => x"c01ec04b",
   129 => x"c1c1f0ff",
   130 => x"87d4fc49",
   131 => x"987086c4",
   132 => x"ff87ca05",
   133 => x"ffc348d4",
   134 => x"cb48c178",
   135 => x"87f1fd87",
   136 => x"ff058bc1",
   137 => x"48c087db",
   138 => x"0e87f1fb",
   139 => x"0e5c5b5e",
   140 => x"fd4cd4ff",
   141 => x"eac687db",
   142 => x"f0e1c01e",
   143 => x"fb49c8c1",
   144 => x"86c487de",
   145 => x"c802a8c1",
   146 => x"87eafe87",
   147 => x"e2c148c0",
   148 => x"87dafa87",
   149 => x"ffcf4970",
   150 => x"eac699ff",
   151 => x"87c802a9",
   152 => x"c087d3fe",
   153 => x"87cbc148",
   154 => x"c07cffc3",
   155 => x"f4fc4bf1",
   156 => x"02987087",
   157 => x"c087ebc0",
   158 => x"f0ffc01e",
   159 => x"fa49fac1",
   160 => x"86c487de",
   161 => x"d9059870",
   162 => x"7cffc387",
   163 => x"ffc3496c",
   164 => x"7c7c7c7c",
   165 => x"0299c0c1",
   166 => x"48c187c4",
   167 => x"48c087d5",
   168 => x"abc287d1",
   169 => x"c087c405",
   170 => x"c187c848",
   171 => x"fdfe058b",
   172 => x"f948c087",
   173 => x"731e87e4",
   174 => x"fce4c21e",
   175 => x"c778c148",
   176 => x"48d0ff4b",
   177 => x"c8fb78c2",
   178 => x"48d0ff87",
   179 => x"1ec078c3",
   180 => x"c1d0e5c0",
   181 => x"c7f949c0",
   182 => x"c186c487",
   183 => x"87c105a8",
   184 => x"05abc24b",
   185 => x"48c087c5",
   186 => x"c187f9c0",
   187 => x"d0ff058b",
   188 => x"87f7fc87",
   189 => x"58c0e5c2",
   190 => x"cd059870",
   191 => x"c01ec187",
   192 => x"d0c1f0ff",
   193 => x"87d8f849",
   194 => x"d4ff86c4",
   195 => x"78ffc348",
   196 => x"c287fcc2",
   197 => x"ff58c4e5",
   198 => x"78c248d0",
   199 => x"c348d4ff",
   200 => x"48c178ff",
   201 => x"0e87f5f7",
   202 => x"5d5c5b5e",
   203 => x"c04b710e",
   204 => x"cdeec54c",
   205 => x"d4ff4adf",
   206 => x"78ffc348",
   207 => x"fec34968",
   208 => x"fdc005a9",
   209 => x"734d7087",
   210 => x"87cc029b",
   211 => x"731e66d0",
   212 => x"87f1f549",
   213 => x"87d686c4",
   214 => x"c448d0ff",
   215 => x"ffc378d1",
   216 => x"4866d07d",
   217 => x"a6d488c1",
   218 => x"05987058",
   219 => x"d4ff87f0",
   220 => x"78ffc348",
   221 => x"059b7378",
   222 => x"d0ff87c5",
   223 => x"c178d048",
   224 => x"8ac14c4a",
   225 => x"87eefe05",
   226 => x"cbf64874",
   227 => x"1e731e87",
   228 => x"4bc04a71",
   229 => x"c348d4ff",
   230 => x"d0ff78ff",
   231 => x"78c3c448",
   232 => x"c348d4ff",
   233 => x"1e7278ff",
   234 => x"c1f0ffc0",
   235 => x"eff549d1",
   236 => x"7086c487",
   237 => x"87d20598",
   238 => x"cc1ec0c8",
   239 => x"e6fd4966",
   240 => x"7086c487",
   241 => x"48d0ff4b",
   242 => x"487378c2",
   243 => x"0e87cdf5",
   244 => x"5d5c5b5e",
   245 => x"c01ec00e",
   246 => x"c9c1f0ff",
   247 => x"87c0f549",
   248 => x"e5c21ed2",
   249 => x"fefc49c4",
   250 => x"c086c887",
   251 => x"d284c14c",
   252 => x"f804acb7",
   253 => x"c4e5c287",
   254 => x"c349bf97",
   255 => x"c0c199c0",
   256 => x"e7c005a9",
   257 => x"cbe5c287",
   258 => x"d049bf97",
   259 => x"cce5c231",
   260 => x"c84abf97",
   261 => x"c2b17232",
   262 => x"bf97cde5",
   263 => x"4c71b14a",
   264 => x"ffffffcf",
   265 => x"ca84c19c",
   266 => x"87e7c134",
   267 => x"97cde5c2",
   268 => x"31c149bf",
   269 => x"e5c299c6",
   270 => x"4abf97ce",
   271 => x"722ab7c7",
   272 => x"c9e5c2b1",
   273 => x"4d4abf97",
   274 => x"e5c29dcf",
   275 => x"4abf97ca",
   276 => x"32ca9ac3",
   277 => x"97cbe5c2",
   278 => x"33c24bbf",
   279 => x"e5c2b273",
   280 => x"4bbf97cc",
   281 => x"c69bc0c3",
   282 => x"b2732bb7",
   283 => x"48c181c2",
   284 => x"49703071",
   285 => x"307548c1",
   286 => x"4c724d70",
   287 => x"947184c1",
   288 => x"adb7c0c8",
   289 => x"c187cc06",
   290 => x"c82db734",
   291 => x"01adb7c0",
   292 => x"7487f4ff",
   293 => x"87c0f248",
   294 => x"5c5b5e0e",
   295 => x"86f80e5d",
   296 => x"48eaedc2",
   297 => x"e5c278c0",
   298 => x"49c01ee2",
   299 => x"c487defb",
   300 => x"05987086",
   301 => x"48c087c5",
   302 => x"c087cec9",
   303 => x"c07ec14d",
   304 => x"49bfd8f5",
   305 => x"4ad8e6c2",
   306 => x"ee4bc871",
   307 => x"987087dc",
   308 => x"c087c205",
   309 => x"d4f5c07e",
   310 => x"e6c249bf",
   311 => x"c8714af4",
   312 => x"87c6ee4b",
   313 => x"c2059870",
   314 => x"6e7ec087",
   315 => x"87fdc002",
   316 => x"bfe8ecc2",
   317 => x"e0edc24d",
   318 => x"487ebf9f",
   319 => x"a8ead6c5",
   320 => x"c287c705",
   321 => x"4dbfe8ec",
   322 => x"486e87ce",
   323 => x"a8d5e9ca",
   324 => x"c087c502",
   325 => x"87f1c748",
   326 => x"1ee2e5c2",
   327 => x"ecf94975",
   328 => x"7086c487",
   329 => x"87c50598",
   330 => x"dcc748c0",
   331 => x"d4f5c087",
   332 => x"e6c249bf",
   333 => x"c8714af4",
   334 => x"87eeec4b",
   335 => x"c8059870",
   336 => x"eaedc287",
   337 => x"da78c148",
   338 => x"d8f5c087",
   339 => x"e6c249bf",
   340 => x"c8714ad8",
   341 => x"87d2ec4b",
   342 => x"c0029870",
   343 => x"48c087c5",
   344 => x"c287e6c6",
   345 => x"bf97e0ed",
   346 => x"a9d5c149",
   347 => x"87cdc005",
   348 => x"97e1edc2",
   349 => x"eac249bf",
   350 => x"c5c002a9",
   351 => x"c648c087",
   352 => x"e5c287c7",
   353 => x"7ebf97e2",
   354 => x"a8e9c348",
   355 => x"87cec002",
   356 => x"ebc3486e",
   357 => x"c5c002a8",
   358 => x"c548c087",
   359 => x"e5c287eb",
   360 => x"49bf97ed",
   361 => x"ccc00599",
   362 => x"eee5c287",
   363 => x"c249bf97",
   364 => x"c5c002a9",
   365 => x"c548c087",
   366 => x"e5c287cf",
   367 => x"48bf97ef",
   368 => x"58e6edc2",
   369 => x"c1484c70",
   370 => x"eaedc288",
   371 => x"f0e5c258",
   372 => x"7549bf97",
   373 => x"f1e5c281",
   374 => x"c84abf97",
   375 => x"7ea17232",
   376 => x"48f7f1c2",
   377 => x"e5c2786e",
   378 => x"48bf97f2",
   379 => x"c258a6c8",
   380 => x"02bfeaed",
   381 => x"c087d4c2",
   382 => x"49bfd4f5",
   383 => x"4af4e6c2",
   384 => x"e94bc871",
   385 => x"987087e4",
   386 => x"87c5c002",
   387 => x"f8c348c0",
   388 => x"e2edc287",
   389 => x"f2c24cbf",
   390 => x"e6c25ccb",
   391 => x"49bf97c7",
   392 => x"e6c231c8",
   393 => x"4abf97c6",
   394 => x"e6c249a1",
   395 => x"4abf97c8",
   396 => x"a17232d0",
   397 => x"c9e6c249",
   398 => x"d84abf97",
   399 => x"49a17232",
   400 => x"c29166c4",
   401 => x"81bff7f1",
   402 => x"59fff1c2",
   403 => x"97cfe6c2",
   404 => x"32c84abf",
   405 => x"97cee6c2",
   406 => x"4aa24bbf",
   407 => x"97d0e6c2",
   408 => x"33d04bbf",
   409 => x"c24aa273",
   410 => x"bf97d1e6",
   411 => x"d89bcf4b",
   412 => x"4aa27333",
   413 => x"5ac3f2c2",
   414 => x"bffff1c2",
   415 => x"748ac24a",
   416 => x"c3f2c292",
   417 => x"78a17248",
   418 => x"c287cac1",
   419 => x"bf97f4e5",
   420 => x"c231c849",
   421 => x"bf97f3e5",
   422 => x"c249a14a",
   423 => x"c259f2ed",
   424 => x"49bfeeed",
   425 => x"ffc731c5",
   426 => x"c229c981",
   427 => x"c259cbf2",
   428 => x"bf97f9e5",
   429 => x"c232c84a",
   430 => x"bf97f8e5",
   431 => x"c44aa24b",
   432 => x"826e9266",
   433 => x"5ac7f2c2",
   434 => x"48fff1c2",
   435 => x"f1c278c0",
   436 => x"a17248fb",
   437 => x"cbf2c278",
   438 => x"fff1c248",
   439 => x"f2c278bf",
   440 => x"f2c248cf",
   441 => x"c278bfc3",
   442 => x"02bfeaed",
   443 => x"7487c9c0",
   444 => x"7030c448",
   445 => x"87c9c07e",
   446 => x"bfc7f2c2",
   447 => x"7030c448",
   448 => x"eeedc27e",
   449 => x"c1786e48",
   450 => x"268ef848",
   451 => x"264c264d",
   452 => x"0e4f264b",
   453 => x"5d5c5b5e",
   454 => x"c24a710e",
   455 => x"02bfeaed",
   456 => x"4b7287cb",
   457 => x"4c722bc7",
   458 => x"c99cffc1",
   459 => x"c84b7287",
   460 => x"c34c722b",
   461 => x"f1c29cff",
   462 => x"c083bff7",
   463 => x"abbfd0f5",
   464 => x"c087d902",
   465 => x"c25bd4f5",
   466 => x"731ee2e5",
   467 => x"87fdf049",
   468 => x"987086c4",
   469 => x"c087c505",
   470 => x"87e6c048",
   471 => x"bfeaedc2",
   472 => x"7487d202",
   473 => x"c291c449",
   474 => x"6981e2e5",
   475 => x"ffffcf4d",
   476 => x"cb9dffff",
   477 => x"c2497487",
   478 => x"e2e5c291",
   479 => x"4d699f81",
   480 => x"c6fe4875",
   481 => x"5b5e0e87",
   482 => x"f80e5d5c",
   483 => x"9c4c7186",
   484 => x"c087c505",
   485 => x"87c1c348",
   486 => x"6e7ea4c8",
   487 => x"d878c048",
   488 => x"87c70266",
   489 => x"bf9766d8",
   490 => x"c087c505",
   491 => x"87e9c248",
   492 => x"49c11ec0",
   493 => x"c487fdce",
   494 => x"9d4d7086",
   495 => x"87c2c102",
   496 => x"4af2edc2",
   497 => x"e24966d8",
   498 => x"987087c5",
   499 => x"87f2c002",
   500 => x"66d84a75",
   501 => x"e24bcb49",
   502 => x"987087ea",
   503 => x"87e2c002",
   504 => x"9d751ec0",
   505 => x"c887c702",
   506 => x"78c048a6",
   507 => x"a6c887c5",
   508 => x"c878c148",
   509 => x"fbcd4966",
   510 => x"7086c487",
   511 => x"fe059d4d",
   512 => x"9d7587fe",
   513 => x"87cfc102",
   514 => x"6e49a5dc",
   515 => x"da786948",
   516 => x"a6c449a5",
   517 => x"78a4c448",
   518 => x"c448699f",
   519 => x"c2780866",
   520 => x"02bfeaed",
   521 => x"a5d487d2",
   522 => x"49699f49",
   523 => x"99ffffc0",
   524 => x"30d04871",
   525 => x"87c27e70",
   526 => x"496e7ec0",
   527 => x"bf66c448",
   528 => x"0866c480",
   529 => x"cc7cc078",
   530 => x"66c449a4",
   531 => x"a4d079bf",
   532 => x"c179c049",
   533 => x"c087c248",
   534 => x"fa8ef848",
   535 => x"5e0e87ed",
   536 => x"0e5d5c5b",
   537 => x"029c4c71",
   538 => x"c887cac1",
   539 => x"026949a4",
   540 => x"d087c2c1",
   541 => x"496c4a66",
   542 => x"5aa6d482",
   543 => x"b94d66d0",
   544 => x"bfe6edc2",
   545 => x"72baff4a",
   546 => x"02997199",
   547 => x"c487e4c0",
   548 => x"496b4ba4",
   549 => x"7087fcf9",
   550 => x"e2edc27b",
   551 => x"816c49bf",
   552 => x"b9757c71",
   553 => x"bfe6edc2",
   554 => x"72baff4a",
   555 => x"05997199",
   556 => x"7587dcff",
   557 => x"87d3f97c",
   558 => x"711e731e",
   559 => x"c7029b4b",
   560 => x"49a3c887",
   561 => x"87c50569",
   562 => x"f7c048c0",
   563 => x"fbf1c287",
   564 => x"a3c44abf",
   565 => x"c2496949",
   566 => x"e2edc289",
   567 => x"a27191bf",
   568 => x"e6edc24a",
   569 => x"996b49bf",
   570 => x"c04aa271",
   571 => x"c85ad4f5",
   572 => x"49721e66",
   573 => x"c487d6ea",
   574 => x"05987086",
   575 => x"48c087c4",
   576 => x"48c187c2",
   577 => x"0e87c8f8",
   578 => x"0e5c5b5e",
   579 => x"d04b711e",
   580 => x"2cc94c66",
   581 => x"c1029b73",
   582 => x"a3c887d4",
   583 => x"c1026949",
   584 => x"edc287cc",
   585 => x"ff49bfe6",
   586 => x"994a6bb9",
   587 => x"03ac717e",
   588 => x"7bc087d1",
   589 => x"c049a3d0",
   590 => x"4aa3cc79",
   591 => x"6a49a3c4",
   592 => x"7287c279",
   593 => x"029c748c",
   594 => x"4987e3c0",
   595 => x"fc49731e",
   596 => x"86c487cc",
   597 => x"c74966d0",
   598 => x"cb0299ff",
   599 => x"e2e5c287",
   600 => x"fd49731e",
   601 => x"86c487d2",
   602 => x"d049a3d0",
   603 => x"f6267966",
   604 => x"5e0e87db",
   605 => x"0e5d5c5b",
   606 => x"a6d086f0",
   607 => x"66e4c059",
   608 => x"0266cc4b",
   609 => x"c84887ca",
   610 => x"6e7e7080",
   611 => x"87c505bf",
   612 => x"ecc348c0",
   613 => x"4c66cc87",
   614 => x"497384d0",
   615 => x"6c48a6c4",
   616 => x"8166c478",
   617 => x"bf6e80c4",
   618 => x"a966c878",
   619 => x"4987c606",
   620 => x"718966c4",
   621 => x"abb7c04b",
   622 => x"4887c401",
   623 => x"c487c2c3",
   624 => x"ffc74866",
   625 => x"6e7e7098",
   626 => x"87c9c102",
   627 => x"6e49c0c8",
   628 => x"c24a7189",
   629 => x"6e4de2e5",
   630 => x"aab77385",
   631 => x"4a87c106",
   632 => x"c4484972",
   633 => x"7c708066",
   634 => x"c1498b72",
   635 => x"0299718a",
   636 => x"e0c087d9",
   637 => x"50154866",
   638 => x"4866e0c0",
   639 => x"e4c080c1",
   640 => x"497258a6",
   641 => x"99718ac1",
   642 => x"c187e705",
   643 => x"4966d01e",
   644 => x"c487cbf9",
   645 => x"abb7c086",
   646 => x"87e3c106",
   647 => x"4d66e0c0",
   648 => x"abb7ffc7",
   649 => x"87e2c006",
   650 => x"66d01e75",
   651 => x"87c8fa49",
   652 => x"6c85c0c8",
   653 => x"80c0c848",
   654 => x"c0c87c70",
   655 => x"d41ec18b",
   656 => x"d9f84966",
   657 => x"c086c887",
   658 => x"e5c287ee",
   659 => x"66d01ee2",
   660 => x"87e4f949",
   661 => x"e5c286c4",
   662 => x"49734ae2",
   663 => x"70806c48",
   664 => x"c149737c",
   665 => x"0299718b",
   666 => x"971287ce",
   667 => x"7385c17d",
   668 => x"718bc149",
   669 => x"87f20599",
   670 => x"01abb7c0",
   671 => x"c187e1fe",
   672 => x"f28ef048",
   673 => x"5e0e87c5",
   674 => x"0e5d5c5b",
   675 => x"029b4b71",
   676 => x"a3c887c7",
   677 => x"c5056d4d",
   678 => x"c048ff87",
   679 => x"a3d087fd",
   680 => x"c7496c4c",
   681 => x"d80599ff",
   682 => x"c9026c87",
   683 => x"731ec187",
   684 => x"87eaf649",
   685 => x"e5c286c4",
   686 => x"49731ee2",
   687 => x"c487f9f7",
   688 => x"6d4a6c86",
   689 => x"87c404aa",
   690 => x"87cf48ff",
   691 => x"727ca2c1",
   692 => x"99ffc749",
   693 => x"81e2e5c2",
   694 => x"f0486997",
   695 => x"731e87ed",
   696 => x"9b4b711e",
   697 => x"87e4c002",
   698 => x"5bcff2c2",
   699 => x"8ac24a73",
   700 => x"bfe2edc2",
   701 => x"f1c29249",
   702 => x"7248bffb",
   703 => x"d3f2c280",
   704 => x"c4487158",
   705 => x"f2edc230",
   706 => x"87edc058",
   707 => x"48cbf2c2",
   708 => x"bffff1c2",
   709 => x"cff2c278",
   710 => x"c3f2c248",
   711 => x"edc278bf",
   712 => x"c902bfea",
   713 => x"e2edc287",
   714 => x"31c449bf",
   715 => x"f2c287c7",
   716 => x"c449bfc7",
   717 => x"f2edc231",
   718 => x"87d3ef59",
   719 => x"5c5b5e0e",
   720 => x"c04a710e",
   721 => x"029a724b",
   722 => x"da87e1c0",
   723 => x"699f49a2",
   724 => x"eaedc24b",
   725 => x"87cf02bf",
   726 => x"9f49a2d4",
   727 => x"c04c4969",
   728 => x"d09cffff",
   729 => x"c087c234",
   730 => x"b349744c",
   731 => x"edfd4973",
   732 => x"87d9ee87",
   733 => x"5c5b5e0e",
   734 => x"86f40e5d",
   735 => x"7ec04a71",
   736 => x"d8029a72",
   737 => x"dee5c287",
   738 => x"c278c048",
   739 => x"c248d6e5",
   740 => x"78bfcff2",
   741 => x"48dae5c2",
   742 => x"bfcbf2c2",
   743 => x"ffedc278",
   744 => x"c250c048",
   745 => x"49bfeeed",
   746 => x"bfdee5c2",
   747 => x"03aa714a",
   748 => x"7287cac4",
   749 => x"0599cf49",
   750 => x"c087eac0",
   751 => x"c248d0f5",
   752 => x"78bfd6e5",
   753 => x"1ee2e5c2",
   754 => x"bfd6e5c2",
   755 => x"d6e5c249",
   756 => x"78a1c148",
   757 => x"f4deff71",
   758 => x"c086c487",
   759 => x"c248ccf5",
   760 => x"cc78e2e5",
   761 => x"ccf5c087",
   762 => x"e0c048bf",
   763 => x"d0f5c080",
   764 => x"dee5c258",
   765 => x"80c148bf",
   766 => x"58e2e5c2",
   767 => x"000d4c27",
   768 => x"bf97bf00",
   769 => x"c2029d4d",
   770 => x"e5c387e3",
   771 => x"dcc202ad",
   772 => x"ccf5c087",
   773 => x"a3cb4bbf",
   774 => x"cf4c1149",
   775 => x"d2c105ac",
   776 => x"df497587",
   777 => x"cd89c199",
   778 => x"f2edc291",
   779 => x"4aa3c181",
   780 => x"a3c35112",
   781 => x"c551124a",
   782 => x"51124aa3",
   783 => x"124aa3c7",
   784 => x"4aa3c951",
   785 => x"a3ce5112",
   786 => x"d051124a",
   787 => x"51124aa3",
   788 => x"124aa3d2",
   789 => x"4aa3d451",
   790 => x"a3d65112",
   791 => x"d851124a",
   792 => x"51124aa3",
   793 => x"124aa3dc",
   794 => x"4aa3de51",
   795 => x"7ec15112",
   796 => x"7487fac0",
   797 => x"0599c849",
   798 => x"7487ebc0",
   799 => x"0599d049",
   800 => x"66dc87d1",
   801 => x"87cbc002",
   802 => x"66dc4973",
   803 => x"0298700f",
   804 => x"6e87d3c0",
   805 => x"87c6c005",
   806 => x"48f2edc2",
   807 => x"f5c050c0",
   808 => x"c248bfcc",
   809 => x"edc287e1",
   810 => x"50c048ff",
   811 => x"eeedc27e",
   812 => x"e5c249bf",
   813 => x"714abfde",
   814 => x"f6fb04aa",
   815 => x"cff2c287",
   816 => x"c8c005bf",
   817 => x"eaedc287",
   818 => x"f8c102bf",
   819 => x"dae5c287",
   820 => x"fee849bf",
   821 => x"c2497087",
   822 => x"c459dee5",
   823 => x"e5c248a6",
   824 => x"c278bfda",
   825 => x"02bfeaed",
   826 => x"c487d8c0",
   827 => x"ffcf4966",
   828 => x"99f8ffff",
   829 => x"c5c002a9",
   830 => x"c04cc087",
   831 => x"4cc187e1",
   832 => x"c487dcc0",
   833 => x"ffcf4966",
   834 => x"02a999f8",
   835 => x"c887c8c0",
   836 => x"78c048a6",
   837 => x"c887c5c0",
   838 => x"78c148a6",
   839 => x"744c66c8",
   840 => x"e0c0059c",
   841 => x"4966c487",
   842 => x"edc289c2",
   843 => x"914abfe2",
   844 => x"bffbf1c2",
   845 => x"d6e5c24a",
   846 => x"78a17248",
   847 => x"48dee5c2",
   848 => x"def978c0",
   849 => x"f448c087",
   850 => x"87ffe68e",
   851 => x"00000000",
   852 => x"ffffffff",
   853 => x"00000d5c",
   854 => x"00000d65",
   855 => x"33544146",
   856 => x"20202032",
   857 => x"54414600",
   858 => x"20203631",
   859 => x"c21e0020",
   860 => x"48bfd4f2",
   861 => x"c905a8dd",
   862 => x"dac2c187",
   863 => x"4a497087",
   864 => x"d4ff87c8",
   865 => x"78ffc348",
   866 => x"48724a68",
   867 => x"c21e4f26",
   868 => x"48bfd4f2",
   869 => x"c605a8dd",
   870 => x"e6c1c187",
   871 => x"ff87d987",
   872 => x"ffc348d4",
   873 => x"48d0ff78",
   874 => x"ff78e1c0",
   875 => x"78d448d4",
   876 => x"48d3f2c2",
   877 => x"50bfd4ff",
   878 => x"ff1e4f26",
   879 => x"e0c048d0",
   880 => x"1e4f2678",
   881 => x"7087e7fe",
   882 => x"c6029949",
   883 => x"a9fbc087",
   884 => x"7187f105",
   885 => x"0e4f2648",
   886 => x"0e5c5b5e",
   887 => x"4cc04b71",
   888 => x"7087cbfe",
   889 => x"c0029949",
   890 => x"ecc087f9",
   891 => x"f2c002a9",
   892 => x"a9fbc087",
   893 => x"87ebc002",
   894 => x"acb766cc",
   895 => x"d087c703",
   896 => x"87c20266",
   897 => x"99715371",
   898 => x"c187c202",
   899 => x"87defd84",
   900 => x"02994970",
   901 => x"ecc087cd",
   902 => x"87c702a9",
   903 => x"05a9fbc0",
   904 => x"d087d5ff",
   905 => x"87c30266",
   906 => x"c07b97c0",
   907 => x"c405a9ec",
   908 => x"c54a7487",
   909 => x"c04a7487",
   910 => x"48728a0a",
   911 => x"4d2687c2",
   912 => x"4b264c26",
   913 => x"fc1e4f26",
   914 => x"497087e4",
   915 => x"aaf0c04a",
   916 => x"c087c904",
   917 => x"c301aaf9",
   918 => x"8af0c087",
   919 => x"04aac1c1",
   920 => x"dac187c9",
   921 => x"87c301aa",
   922 => x"728af7c0",
   923 => x"0e4f2648",
   924 => x"0e5c5b5e",
   925 => x"d4ff4a71",
   926 => x"c049724c",
   927 => x"4b7087e9",
   928 => x"87c2029b",
   929 => x"d0ff8bc1",
   930 => x"c178c548",
   931 => x"49737cd5",
   932 => x"e7c131c6",
   933 => x"4abf97c9",
   934 => x"70b07148",
   935 => x"48d0ff7c",
   936 => x"487378c4",
   937 => x"0e87d9fe",
   938 => x"5d5c5b5e",
   939 => x"7186f40e",
   940 => x"48a6c44c",
   941 => x"a4c878c0",
   942 => x"bf976e7e",
   943 => x"a9c1c149",
   944 => x"c987dd05",
   945 => x"699749a4",
   946 => x"a9d2c149",
   947 => x"ca87d105",
   948 => x"699749a4",
   949 => x"a9c3c149",
   950 => x"df87c505",
   951 => x"87e1c248",
   952 => x"c087ebfa",
   953 => x"c6fec04b",
   954 => x"c049bf97",
   955 => x"87cf04a9",
   956 => x"c187d0fb",
   957 => x"c6fec083",
   958 => x"ab49bf97",
   959 => x"c087f106",
   960 => x"bf97c6fe",
   961 => x"f987cf02",
   962 => x"497087e4",
   963 => x"87c60299",
   964 => x"05a9ecc0",
   965 => x"4bc087f1",
   966 => x"7087d3f9",
   967 => x"87cef94d",
   968 => x"f958a6cc",
   969 => x"4a7087c8",
   970 => x"976e83c1",
   971 => x"02ad49bf",
   972 => x"ffc087c7",
   973 => x"eac005ad",
   974 => x"49a4c987",
   975 => x"c8496997",
   976 => x"c702a966",
   977 => x"ffc04887",
   978 => x"87d705a8",
   979 => x"9749a4ca",
   980 => x"02aa4969",
   981 => x"ffc087c6",
   982 => x"87c705aa",
   983 => x"c148a6c4",
   984 => x"c087d378",
   985 => x"c602adec",
   986 => x"adfbc087",
   987 => x"c087c705",
   988 => x"48a6c44b",
   989 => x"66c478c1",
   990 => x"87dcfe02",
   991 => x"7387fbf8",
   992 => x"fa8ef448",
   993 => x"0e0087f8",
   994 => x"5d5c5b5e",
   995 => x"7186f80e",
   996 => x"4bd4ff4d",
   997 => x"f2c21e75",
   998 => x"dfff49d8",
   999 => x"86c487e7",
  1000 => x"c4029870",
  1001 => x"e7c187fb",
  1002 => x"757ebfcb",
  1003 => x"87fffa49",
  1004 => x"c005a8de",
  1005 => x"497587eb",
  1006 => x"87f9f6c0",
  1007 => x"db029870",
  1008 => x"fcf6c287",
  1009 => x"e1c01ebf",
  1010 => x"c8f4c049",
  1011 => x"c186c487",
  1012 => x"c048c9e7",
  1013 => x"c8f7c250",
  1014 => x"87ebfe49",
  1015 => x"c2c448c1",
  1016 => x"48d0ff87",
  1017 => x"d6c178c5",
  1018 => x"754ac07b",
  1019 => x"7b1149a2",
  1020 => x"b7cb82c1",
  1021 => x"87f304aa",
  1022 => x"ffc34acc",
  1023 => x"c082c17b",
  1024 => x"04aab7e0",
  1025 => x"d0ff87f4",
  1026 => x"c378c448",
  1027 => x"78c57bff",
  1028 => x"c17bd3c1",
  1029 => x"6e78c47b",
  1030 => x"a8b7c048",
  1031 => x"87f0c206",
  1032 => x"bfe0f2c2",
  1033 => x"74486e4c",
  1034 => x"747e7088",
  1035 => x"fdc1029c",
  1036 => x"e2e5c287",
  1037 => x"48a6c44d",
  1038 => x"8c78c0c8",
  1039 => x"03acb7c0",
  1040 => x"c0c887c6",
  1041 => x"4cc078a4",
  1042 => x"97d3f2c2",
  1043 => x"99d049bf",
  1044 => x"c087d102",
  1045 => x"d8f2c21e",
  1046 => x"87dce149",
  1047 => x"497086c4",
  1048 => x"87eec04a",
  1049 => x"1ee2e5c2",
  1050 => x"49d8f2c2",
  1051 => x"c487c9e1",
  1052 => x"4a497086",
  1053 => x"c848d0ff",
  1054 => x"d4c178c5",
  1055 => x"c47b157b",
  1056 => x"88c14866",
  1057 => x"7058a6c8",
  1058 => x"f0ff0598",
  1059 => x"48d0ff87",
  1060 => x"9a7278c4",
  1061 => x"c087c505",
  1062 => x"87c7c148",
  1063 => x"f2c21ec1",
  1064 => x"deff49d8",
  1065 => x"86c487f8",
  1066 => x"fe059c74",
  1067 => x"486e87c3",
  1068 => x"06a8b7c0",
  1069 => x"f2c287d1",
  1070 => x"78c048d8",
  1071 => x"78c080d0",
  1072 => x"f2c280f4",
  1073 => x"6e78bfe4",
  1074 => x"a8b7c048",
  1075 => x"87d0fd01",
  1076 => x"c548d0ff",
  1077 => x"7bd3c178",
  1078 => x"78c47bc0",
  1079 => x"c2c048c1",
  1080 => x"f848c087",
  1081 => x"264d268e",
  1082 => x"264b264c",
  1083 => x"5b5e0e4f",
  1084 => x"1e0e5d5c",
  1085 => x"4cc04b71",
  1086 => x"c004ab4d",
  1087 => x"fac087e8",
  1088 => x"9d751ee7",
  1089 => x"c087c402",
  1090 => x"c187c24a",
  1091 => x"e949724a",
  1092 => x"86c487e2",
  1093 => x"84c17e70",
  1094 => x"87c2056e",
  1095 => x"85c14c73",
  1096 => x"ff06ac73",
  1097 => x"486e87d8",
  1098 => x"87f9fe26",
  1099 => x"c44a711e",
  1100 => x"87c50566",
  1101 => x"cef94972",
  1102 => x"0e4f2687",
  1103 => x"5d5c5b5e",
  1104 => x"4c711e0e",
  1105 => x"c291de49",
  1106 => x"714dc0f3",
  1107 => x"026d9785",
  1108 => x"c287dcc1",
  1109 => x"4abfecf2",
  1110 => x"49728274",
  1111 => x"7087cefe",
  1112 => x"c0026e7e",
  1113 => x"f2c287f2",
  1114 => x"4a6e4bf4",
  1115 => x"fcfe49cb",
  1116 => x"4b7487f6",
  1117 => x"e7c193cb",
  1118 => x"83c483dd",
  1119 => x"7bf3c6c1",
  1120 => x"cbc14974",
  1121 => x"7b7587d0",
  1122 => x"97cae7c1",
  1123 => x"c21e49bf",
  1124 => x"fe49f4f2",
  1125 => x"86c487d6",
  1126 => x"cac14974",
  1127 => x"49c087f8",
  1128 => x"87d7ccc1",
  1129 => x"48d4f2c2",
  1130 => x"49c178c0",
  1131 => x"2687d9dd",
  1132 => x"4c87f2fc",
  1133 => x"6964616f",
  1134 => x"2e2e676e",
  1135 => x"5e0e002e",
  1136 => x"710e5c5b",
  1137 => x"f2c24a4b",
  1138 => x"7282bfec",
  1139 => x"87ddfc49",
  1140 => x"029c4c70",
  1141 => x"e54987c4",
  1142 => x"f2c287e2",
  1143 => x"78c048ec",
  1144 => x"e3dc49c1",
  1145 => x"87fffb87",
  1146 => x"5c5b5e0e",
  1147 => x"86f40e5d",
  1148 => x"4de2e5c2",
  1149 => x"a6c44cc0",
  1150 => x"c278c048",
  1151 => x"49bfecf2",
  1152 => x"c106a9c0",
  1153 => x"e5c287c1",
  1154 => x"029848e2",
  1155 => x"c087f8c0",
  1156 => x"c81ee7fa",
  1157 => x"87c70266",
  1158 => x"c048a6c4",
  1159 => x"c487c578",
  1160 => x"78c148a6",
  1161 => x"e54966c4",
  1162 => x"86c487ca",
  1163 => x"84c14d70",
  1164 => x"c14866c4",
  1165 => x"58a6c880",
  1166 => x"bfecf2c2",
  1167 => x"c603ac49",
  1168 => x"059d7587",
  1169 => x"c087c8ff",
  1170 => x"029d754c",
  1171 => x"c087e0c3",
  1172 => x"c81ee7fa",
  1173 => x"87c70266",
  1174 => x"c048a6cc",
  1175 => x"cc87c578",
  1176 => x"78c148a6",
  1177 => x"e44966cc",
  1178 => x"86c487ca",
  1179 => x"026e7e70",
  1180 => x"6e87e9c2",
  1181 => x"9781cb49",
  1182 => x"99d04969",
  1183 => x"87d6c102",
  1184 => x"4afec6c1",
  1185 => x"91cb4974",
  1186 => x"81dde7c1",
  1187 => x"81c87972",
  1188 => x"7451ffc3",
  1189 => x"c291de49",
  1190 => x"714dc0f3",
  1191 => x"97c1c285",
  1192 => x"49a5c17d",
  1193 => x"c251e0c0",
  1194 => x"bf97f2ed",
  1195 => x"c187d202",
  1196 => x"4ba5c284",
  1197 => x"4af2edc2",
  1198 => x"f7fe49db",
  1199 => x"dbc187ea",
  1200 => x"49a5cd87",
  1201 => x"84c151c0",
  1202 => x"6e4ba5c2",
  1203 => x"fe49cb4a",
  1204 => x"c187d5f7",
  1205 => x"c4c187c6",
  1206 => x"49744afb",
  1207 => x"e7c191cb",
  1208 => x"797281dd",
  1209 => x"97f2edc2",
  1210 => x"87d802bf",
  1211 => x"91de4974",
  1212 => x"f3c284c1",
  1213 => x"83714bc0",
  1214 => x"4af2edc2",
  1215 => x"f6fe49dd",
  1216 => x"87d887e6",
  1217 => x"93de4b74",
  1218 => x"83c0f3c2",
  1219 => x"c049a3cb",
  1220 => x"7384c151",
  1221 => x"49cb4a6e",
  1222 => x"87ccf6fe",
  1223 => x"c14866c4",
  1224 => x"58a6c880",
  1225 => x"c003acc7",
  1226 => x"056e87c5",
  1227 => x"7487e0fc",
  1228 => x"f68ef448",
  1229 => x"731e87ef",
  1230 => x"494b711e",
  1231 => x"e7c191cb",
  1232 => x"a1c881dd",
  1233 => x"c9e7c14a",
  1234 => x"c9501248",
  1235 => x"fec04aa1",
  1236 => x"501248c6",
  1237 => x"e7c181ca",
  1238 => x"501148ca",
  1239 => x"97cae7c1",
  1240 => x"c01e49bf",
  1241 => x"87c4f749",
  1242 => x"48d4f2c2",
  1243 => x"49c178de",
  1244 => x"2687d5d6",
  1245 => x"1e87f2f5",
  1246 => x"cb494a71",
  1247 => x"dde7c191",
  1248 => x"1181c881",
  1249 => x"d8f2c248",
  1250 => x"ecf2c258",
  1251 => x"c178c048",
  1252 => x"87f4d549",
  1253 => x"c01e4f26",
  1254 => x"dec4c149",
  1255 => x"1e4f2687",
  1256 => x"d2029971",
  1257 => x"f2e8c187",
  1258 => x"f750c048",
  1259 => x"f7cdc180",
  1260 => x"d6e7c140",
  1261 => x"c187ce78",
  1262 => x"c148eee8",
  1263 => x"fc78cfe7",
  1264 => x"d6cec180",
  1265 => x"0e4f2678",
  1266 => x"0e5c5b5e",
  1267 => x"cb4a4c71",
  1268 => x"dde7c192",
  1269 => x"49a2c882",
  1270 => x"974ba2c9",
  1271 => x"971e4b6b",
  1272 => x"ca1e4969",
  1273 => x"c0491282",
  1274 => x"c087cae5",
  1275 => x"87d8d449",
  1276 => x"c1c14974",
  1277 => x"8ef887e0",
  1278 => x"1e87ecf3",
  1279 => x"4b711e73",
  1280 => x"87c3ff49",
  1281 => x"fefe4973",
  1282 => x"87ddf387",
  1283 => x"711e731e",
  1284 => x"4aa3c64b",
  1285 => x"c187db02",
  1286 => x"87d6028a",
  1287 => x"dac1028a",
  1288 => x"c0028a87",
  1289 => x"028a87fc",
  1290 => x"8a87e1c0",
  1291 => x"c187cb02",
  1292 => x"49c787db",
  1293 => x"c187c0fd",
  1294 => x"f2c287de",
  1295 => x"c102bfec",
  1296 => x"c14887cb",
  1297 => x"f0f2c288",
  1298 => x"87c1c158",
  1299 => x"bff0f2c2",
  1300 => x"87f9c002",
  1301 => x"bfecf2c2",
  1302 => x"c280c148",
  1303 => x"c058f0f2",
  1304 => x"f2c287eb",
  1305 => x"c649bfec",
  1306 => x"f0f2c289",
  1307 => x"a9b7c059",
  1308 => x"c287da03",
  1309 => x"c048ecf2",
  1310 => x"c287d278",
  1311 => x"02bff0f2",
  1312 => x"f2c287cb",
  1313 => x"c648bfec",
  1314 => x"f0f2c280",
  1315 => x"d149c058",
  1316 => x"497387f6",
  1317 => x"87fefec0",
  1318 => x"1e87cef1",
  1319 => x"4b711e73",
  1320 => x"48d4f2c2",
  1321 => x"49c078dd",
  1322 => x"7387ddd1",
  1323 => x"e5fec049",
  1324 => x"87f5f087",
  1325 => x"5c5b5e0e",
  1326 => x"ccff0e5d",
  1327 => x"59a6d886",
  1328 => x"c048a6c8",
  1329 => x"c180c478",
  1330 => x"c47866c8",
  1331 => x"c278c180",
  1332 => x"c148f0f2",
  1333 => x"d4f2c278",
  1334 => x"a8de48bf",
  1335 => x"f487cb05",
  1336 => x"497087c6",
  1337 => x"cf59a6cc",
  1338 => x"e1e287d0",
  1339 => x"87d3e387",
  1340 => x"7087fbe1",
  1341 => x"0566d44c",
  1342 => x"c187fcc1",
  1343 => x"c44866c4",
  1344 => x"c47e7080",
  1345 => x"bf6e48a6",
  1346 => x"c11e7278",
  1347 => x"c848efe3",
  1348 => x"a1c84966",
  1349 => x"7141204a",
  1350 => x"87f905aa",
  1351 => x"4a265110",
  1352 => x"4866c4c1",
  1353 => x"78f6ccc1",
  1354 => x"c749bf6e",
  1355 => x"c1517481",
  1356 => x"c84966c4",
  1357 => x"c151c181",
  1358 => x"c94966c4",
  1359 => x"c151c081",
  1360 => x"ca4966c4",
  1361 => x"c051c081",
  1362 => x"cf02acfb",
  1363 => x"d81ec187",
  1364 => x"bf66c81e",
  1365 => x"e181c849",
  1366 => x"86c887fd",
  1367 => x"4866c8c1",
  1368 => x"c701a8c0",
  1369 => x"48a6c887",
  1370 => x"87ce78c1",
  1371 => x"4866c8c1",
  1372 => x"a6d088c1",
  1373 => x"e187c358",
  1374 => x"a6d887c9",
  1375 => x"7478c248",
  1376 => x"f1cc029c",
  1377 => x"4866c887",
  1378 => x"a866ccc1",
  1379 => x"87e6cc03",
  1380 => x"c048a6dc",
  1381 => x"c080c478",
  1382 => x"d1dfff78",
  1383 => x"d44c7087",
  1384 => x"a8dd4866",
  1385 => x"c087c705",
  1386 => x"d448a6e0",
  1387 => x"d0c17866",
  1388 => x"ebc005ac",
  1389 => x"f5deff87",
  1390 => x"f1deff87",
  1391 => x"c04c7087",
  1392 => x"c605acec",
  1393 => x"fadfff87",
  1394 => x"c14c7087",
  1395 => x"c805acd0",
  1396 => x"4866d087",
  1397 => x"a6d480c1",
  1398 => x"acd0c158",
  1399 => x"87d5ff02",
  1400 => x"48a6e4c0",
  1401 => x"c07866d4",
  1402 => x"c04866e0",
  1403 => x"05a866e4",
  1404 => x"c087d5ca",
  1405 => x"c048a6e8",
  1406 => x"80dcff78",
  1407 => x"4d7478c0",
  1408 => x"028dfbc0",
  1409 => x"c987dbc9",
  1410 => x"87db028d",
  1411 => x"c1028dc2",
  1412 => x"8dc987f7",
  1413 => x"87d8c402",
  1414 => x"c1028dc4",
  1415 => x"8dc187c1",
  1416 => x"87ccc402",
  1417 => x"c887f5c8",
  1418 => x"91cb4966",
  1419 => x"8166c4c1",
  1420 => x"6a4aa1c4",
  1421 => x"c11e717e",
  1422 => x"c448fbe3",
  1423 => x"a1cc4966",
  1424 => x"7141204a",
  1425 => x"f8ff05aa",
  1426 => x"26511087",
  1427 => x"dbd2c149",
  1428 => x"d9dcff79",
  1429 => x"c44c7087",
  1430 => x"78c148a6",
  1431 => x"dc87c3c8",
  1432 => x"f0c048a6",
  1433 => x"c5dcff78",
  1434 => x"c04c7087",
  1435 => x"c002acec",
  1436 => x"e0c087c4",
  1437 => x"ecc05ca6",
  1438 => x"87cd02ac",
  1439 => x"87eedbff",
  1440 => x"ecc04c70",
  1441 => x"f3ff05ac",
  1442 => x"acecc087",
  1443 => x"87c4c002",
  1444 => x"87dadbff",
  1445 => x"1eca1ec0",
  1446 => x"cb4966d0",
  1447 => x"66ccc191",
  1448 => x"cc807148",
  1449 => x"66c858a6",
  1450 => x"d080c448",
  1451 => x"66cc58a6",
  1452 => x"dcff49bf",
  1453 => x"1ec187e1",
  1454 => x"66d41ede",
  1455 => x"dcff49bf",
  1456 => x"86d087d5",
  1457 => x"09c04970",
  1458 => x"a6f0c089",
  1459 => x"66ecc059",
  1460 => x"06a8c048",
  1461 => x"c087eec0",
  1462 => x"dd4866ec",
  1463 => x"e4c003a8",
  1464 => x"bf66c487",
  1465 => x"66ecc049",
  1466 => x"51e0c081",
  1467 => x"4966ecc0",
  1468 => x"66c481c1",
  1469 => x"c1c281bf",
  1470 => x"66ecc051",
  1471 => x"c481c249",
  1472 => x"c081bf66",
  1473 => x"c1486e51",
  1474 => x"6e78f6cc",
  1475 => x"d881c849",
  1476 => x"496e5166",
  1477 => x"66d081c9",
  1478 => x"ca496e51",
  1479 => x"5166dc81",
  1480 => x"c14866d8",
  1481 => x"58a6dc80",
  1482 => x"c180ec48",
  1483 => x"87f2c478",
  1484 => x"87d2dcff",
  1485 => x"f0c04970",
  1486 => x"dcff59a6",
  1487 => x"497087c8",
  1488 => x"59a6e0c0",
  1489 => x"c04866dc",
  1490 => x"c005a8ec",
  1491 => x"a6dc87ca",
  1492 => x"66ecc048",
  1493 => x"87c4c078",
  1494 => x"87d2d8ff",
  1495 => x"cb4966c8",
  1496 => x"66c4c191",
  1497 => x"70807148",
  1498 => x"c84a6e7e",
  1499 => x"ca496e82",
  1500 => x"66ecc081",
  1501 => x"4966dc51",
  1502 => x"ecc081c1",
  1503 => x"48c18966",
  1504 => x"49703071",
  1505 => x"977189c1",
  1506 => x"dcf6c27a",
  1507 => x"ecc049bf",
  1508 => x"6a972966",
  1509 => x"9871484a",
  1510 => x"58a6f4c0",
  1511 => x"81c4496e",
  1512 => x"786948a6",
  1513 => x"4866e4c0",
  1514 => x"a866e0c0",
  1515 => x"87c8c002",
  1516 => x"c048a6dc",
  1517 => x"87c5c078",
  1518 => x"c148a6dc",
  1519 => x"1e66dc78",
  1520 => x"cc1ee0c0",
  1521 => x"d8ff4966",
  1522 => x"86c887cd",
  1523 => x"b7c04c70",
  1524 => x"dbc106ac",
  1525 => x"4866c487",
  1526 => x"a6c88074",
  1527 => x"49e0c058",
  1528 => x"66c48974",
  1529 => x"f8e3c14b",
  1530 => x"e2fe714a",
  1531 => x"66c487fa",
  1532 => x"c880c248",
  1533 => x"e8c058a6",
  1534 => x"80c14866",
  1535 => x"58a6ecc0",
  1536 => x"4966f0c0",
  1537 => x"a97081c1",
  1538 => x"87c5c002",
  1539 => x"c2c04dc0",
  1540 => x"754dc187",
  1541 => x"49a4c21e",
  1542 => x"7148e0c0",
  1543 => x"1e497088",
  1544 => x"ff4966cc",
  1545 => x"c887f0d6",
  1546 => x"a8b7c086",
  1547 => x"87c6ff01",
  1548 => x"0266e8c0",
  1549 => x"6e87d1c0",
  1550 => x"c081c949",
  1551 => x"6e5166e8",
  1552 => x"c7cfc148",
  1553 => x"87ccc078",
  1554 => x"81c9496e",
  1555 => x"486e51c2",
  1556 => x"78fbcfc1",
  1557 => x"c148a6c4",
  1558 => x"87c6c078",
  1559 => x"87e3d5ff",
  1560 => x"66c44c70",
  1561 => x"87f5c002",
  1562 => x"cc4866c8",
  1563 => x"c004a866",
  1564 => x"66c887cb",
  1565 => x"cc80c148",
  1566 => x"e0c058a6",
  1567 => x"4866cc87",
  1568 => x"a6d088c1",
  1569 => x"87d5c058",
  1570 => x"05acc6c1",
  1571 => x"d887c8c0",
  1572 => x"80c14866",
  1573 => x"ff58a6dc",
  1574 => x"7087e8d4",
  1575 => x"4866d04c",
  1576 => x"a6d480c1",
  1577 => x"029c7458",
  1578 => x"c887cbc0",
  1579 => x"ccc14866",
  1580 => x"f304a866",
  1581 => x"d4ff87da",
  1582 => x"66c887c0",
  1583 => x"03a8c748",
  1584 => x"c287e5c0",
  1585 => x"c048f0f2",
  1586 => x"4966c878",
  1587 => x"c4c191cb",
  1588 => x"a1c48166",
  1589 => x"c04a6a4a",
  1590 => x"66c87952",
  1591 => x"cc80c148",
  1592 => x"a8c758a6",
  1593 => x"87dbff04",
  1594 => x"ff8eccff",
  1595 => x"4c87f6df",
  1596 => x"2064616f",
  1597 => x"00202e2a",
  1598 => x"4400203a",
  1599 => x"53205049",
  1600 => x"63746977",
  1601 => x"00736568",
  1602 => x"711e731e",
  1603 => x"c6029b4b",
  1604 => x"ecf2c287",
  1605 => x"c778c048",
  1606 => x"ecf2c21e",
  1607 => x"c11e49bf",
  1608 => x"c21edde7",
  1609 => x"49bfd4f2",
  1610 => x"cc87c9ee",
  1611 => x"d4f2c286",
  1612 => x"eae949bf",
  1613 => x"029b7387",
  1614 => x"e7c187c8",
  1615 => x"edc049dd",
  1616 => x"deff87e6",
  1617 => x"c71e87e3",
  1618 => x"49c187cd",
  1619 => x"fe87f9fe",
  1620 => x"7087e3e5",
  1621 => x"87cd0298",
  1622 => x"87fcecfe",
  1623 => x"c4029870",
  1624 => x"c24ac187",
  1625 => x"724ac087",
  1626 => x"87ce059a",
  1627 => x"e6c11ec0",
  1628 => x"f9c049db",
  1629 => x"86c487d0",
  1630 => x"fbc087fe",
  1631 => x"1ec087f3",
  1632 => x"49e6e6c1",
  1633 => x"87fef8c0",
  1634 => x"fdc01ec0",
  1635 => x"497087f9",
  1636 => x"87f2f8c0",
  1637 => x"f887ffc2",
  1638 => x"534f268e",
  1639 => x"61662044",
  1640 => x"64656c69",
  1641 => x"6f42002e",
  1642 => x"6e69746f",
  1643 => x"2e2e2e67",
  1644 => x"f2c21e00",
  1645 => x"78c048ec",
  1646 => x"48d4f2c2",
  1647 => x"c5fe78c0",
  1648 => x"e1fdc087",
  1649 => x"2648c087",
  1650 => x"0100004f",
  1651 => x"80000000",
  1652 => x"69784520",
  1653 => x"20800074",
  1654 => x"6b636142",
  1655 => x"00137700",
  1656 => x"002cc000",
  1657 => x"00000000",
  1658 => x"00001377",
  1659 => x"00002cde",
  1660 => x"77000000",
  1661 => x"fc000013",
  1662 => x"0000002c",
  1663 => x"13770000",
  1664 => x"2d1a0000",
  1665 => x"00000000",
  1666 => x"00137700",
  1667 => x"002d3800",
  1668 => x"00000000",
  1669 => x"00001377",
  1670 => x"00002d56",
  1671 => x"77000000",
  1672 => x"74000013",
  1673 => x"0000002d",
  1674 => x"13770000",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"00140c00",
  1678 => x"00000000",
  1679 => x"00000000",
  1680 => x"48f0fe1e",
  1681 => x"09cd78c0",
  1682 => x"4f260979",
  1683 => x"f0fe1e1e",
  1684 => x"26487ebf",
  1685 => x"fe1e4f26",
  1686 => x"78c148f0",
  1687 => x"fe1e4f26",
  1688 => x"78c048f0",
  1689 => x"711e4f26",
  1690 => x"5252c04a",
  1691 => x"5e0e4f26",
  1692 => x"0e5d5c5b",
  1693 => x"4d7186f4",
  1694 => x"c17e6d97",
  1695 => x"6c974ca5",
  1696 => x"58a6c848",
  1697 => x"66c4486e",
  1698 => x"87c505a8",
  1699 => x"e6c048ff",
  1700 => x"87caff87",
  1701 => x"9749a5c2",
  1702 => x"a3714b6c",
  1703 => x"4b6b974b",
  1704 => x"6e7e6c97",
  1705 => x"c880c148",
  1706 => x"98c758a6",
  1707 => x"7058a6cc",
  1708 => x"e1fe7c97",
  1709 => x"f4487387",
  1710 => x"264d268e",
  1711 => x"264b264c",
  1712 => x"5b5e0e4f",
  1713 => x"86f40e5c",
  1714 => x"66d84c71",
  1715 => x"9affc34a",
  1716 => x"974ba4c2",
  1717 => x"a173496c",
  1718 => x"97517249",
  1719 => x"486e7e6c",
  1720 => x"a6c880c1",
  1721 => x"cc98c758",
  1722 => x"547058a6",
  1723 => x"caff8ef4",
  1724 => x"fd1e1e87",
  1725 => x"bfe087e8",
  1726 => x"e0c0494a",
  1727 => x"cb0299c0",
  1728 => x"c21e7287",
  1729 => x"fe49d2f6",
  1730 => x"86c487f7",
  1731 => x"7087fdfc",
  1732 => x"87c2fd7e",
  1733 => x"1e4f2626",
  1734 => x"49d2f6c2",
  1735 => x"c187c7fd",
  1736 => x"fc49f1eb",
  1737 => x"c7c487da",
  1738 => x"1e4f2687",
  1739 => x"c848d0ff",
  1740 => x"d4ff78e1",
  1741 => x"c478c548",
  1742 => x"87c30266",
  1743 => x"c878e0c3",
  1744 => x"87c60266",
  1745 => x"c348d4ff",
  1746 => x"d4ff78f0",
  1747 => x"ff787148",
  1748 => x"e1c848d0",
  1749 => x"78e0c078",
  1750 => x"5e0e4f26",
  1751 => x"710e5c5b",
  1752 => x"d2f6c24c",
  1753 => x"87c6fc49",
  1754 => x"b7c04a70",
  1755 => x"e2c204aa",
  1756 => x"aaf0c387",
  1757 => x"c187c905",
  1758 => x"c148dff0",
  1759 => x"87c3c278",
  1760 => x"05aae0c3",
  1761 => x"f0c187c9",
  1762 => x"78c148e3",
  1763 => x"c187f4c1",
  1764 => x"02bfe3f0",
  1765 => x"c0c287c6",
  1766 => x"87c24ba2",
  1767 => x"9c744b72",
  1768 => x"c187d105",
  1769 => x"1ebfdff0",
  1770 => x"bfe3f0c1",
  1771 => x"fd49721e",
  1772 => x"86c887f9",
  1773 => x"bfdff0c1",
  1774 => x"87e0c002",
  1775 => x"b7c44973",
  1776 => x"f1c19129",
  1777 => x"4a7381ff",
  1778 => x"92c29acf",
  1779 => x"307248c1",
  1780 => x"baff4a70",
  1781 => x"98694872",
  1782 => x"87db7970",
  1783 => x"b7c44973",
  1784 => x"f1c19129",
  1785 => x"4a7381ff",
  1786 => x"92c29acf",
  1787 => x"307248c3",
  1788 => x"69484a70",
  1789 => x"c17970b0",
  1790 => x"c048e3f0",
  1791 => x"dff0c178",
  1792 => x"c278c048",
  1793 => x"f949d2f6",
  1794 => x"4a7087e4",
  1795 => x"03aab7c0",
  1796 => x"c087defd",
  1797 => x"2687c248",
  1798 => x"264c264d",
  1799 => x"004f264b",
  1800 => x"00000000",
  1801 => x"1e000000",
  1802 => x"fc494a71",
  1803 => x"4f2687ec",
  1804 => x"724ac01e",
  1805 => x"c191c449",
  1806 => x"c081fff1",
  1807 => x"d082c179",
  1808 => x"ee04aab7",
  1809 => x"0e4f2687",
  1810 => x"5d5c5b5e",
  1811 => x"f84d710e",
  1812 => x"4a7587cc",
  1813 => x"922ab7c4",
  1814 => x"82fff1c1",
  1815 => x"9ccf4c75",
  1816 => x"496a94c2",
  1817 => x"c32b744b",
  1818 => x"7448c29b",
  1819 => x"ff4c7030",
  1820 => x"714874bc",
  1821 => x"f77a7098",
  1822 => x"487387dc",
  1823 => x"0087d8fe",
  1824 => x"00000000",
  1825 => x"00000000",
  1826 => x"00000000",
  1827 => x"00000000",
  1828 => x"00000000",
  1829 => x"00000000",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00000000",
  1834 => x"00000000",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"1e000000",
  1840 => x"c848d0ff",
  1841 => x"487178e1",
  1842 => x"7808d4ff",
  1843 => x"ff4866c4",
  1844 => x"267808d4",
  1845 => x"4a711e4f",
  1846 => x"1e4966c4",
  1847 => x"deff4972",
  1848 => x"48d0ff87",
  1849 => x"2678e0c0",
  1850 => x"731e4f26",
  1851 => x"c84b711e",
  1852 => x"731e4966",
  1853 => x"a2e0c14a",
  1854 => x"87d9ff49",
  1855 => x"2687c426",
  1856 => x"264c264d",
  1857 => x"1e4f264b",
  1858 => x"c34ad4ff",
  1859 => x"d0ff7aff",
  1860 => x"78e1c048",
  1861 => x"f6c27ade",
  1862 => x"497abfdc",
  1863 => x"7028c848",
  1864 => x"d048717a",
  1865 => x"717a7028",
  1866 => x"7028d848",
  1867 => x"48d0ff7a",
  1868 => x"2678e0c0",
  1869 => x"5b5e0e4f",
  1870 => x"710e5d5c",
  1871 => x"dcf6c24c",
  1872 => x"744b4dbf",
  1873 => x"9b66d02b",
  1874 => x"66d483c1",
  1875 => x"87c204ab",
  1876 => x"4a744bc0",
  1877 => x"724966d0",
  1878 => x"75b9ff31",
  1879 => x"72487399",
  1880 => x"484a7030",
  1881 => x"f6c2b071",
  1882 => x"dafe58e0",
  1883 => x"264d2687",
  1884 => x"264b264c",
  1885 => x"5b5e0e4f",
  1886 => x"1e0e5d5c",
  1887 => x"f6c24c71",
  1888 => x"4ac04be0",
  1889 => x"fe49f4c0",
  1890 => x"7487edcc",
  1891 => x"e0f6c21e",
  1892 => x"f0e7fe49",
  1893 => x"7086c487",
  1894 => x"c0029949",
  1895 => x"1ec487ea",
  1896 => x"c21e4da6",
  1897 => x"fe49e0f6",
  1898 => x"c887c7ef",
  1899 => x"02987086",
  1900 => x"4a7587d6",
  1901 => x"49fef7c1",
  1902 => x"cafe4bc4",
  1903 => x"987087ec",
  1904 => x"c087ca02",
  1905 => x"87edc048",
  1906 => x"e8c048c0",
  1907 => x"87f3c087",
  1908 => x"7087c4c1",
  1909 => x"87c80298",
  1910 => x"7087fcc0",
  1911 => x"87f80598",
  1912 => x"bfc0f7c2",
  1913 => x"c287cc02",
  1914 => x"c248dcf6",
  1915 => x"78bfc0f7",
  1916 => x"c187d4fc",
  1917 => x"4d262648",
  1918 => x"4b264c26",
  1919 => x"415b4f26",
  1920 => x"1e004352",
  1921 => x"f6c21ec0",
  1922 => x"ebfe49e0",
  1923 => x"f6c287f9",
  1924 => x"78c048f8",
  1925 => x"0e4f2626",
  1926 => x"5d5c5b5e",
  1927 => x"c086f40e",
  1928 => x"f8f6c27e",
  1929 => x"b7c348bf",
  1930 => x"87d103a8",
  1931 => x"bff8f6c2",
  1932 => x"c280c148",
  1933 => x"c058fcf6",
  1934 => x"d9c648fb",
  1935 => x"e0f6c287",
  1936 => x"c1f1fe49",
  1937 => x"c04c7087",
  1938 => x"c403acb7",
  1939 => x"c5c64887",
  1940 => x"f8f6c287",
  1941 => x"8ac34abf",
  1942 => x"c187d802",
  1943 => x"c7c5028a",
  1944 => x"c2028a87",
  1945 => x"028a87f2",
  1946 => x"8a87cfc1",
  1947 => x"87dec302",
  1948 => x"c087d9c5",
  1949 => x"5ca6c84d",
  1950 => x"92c44a75",
  1951 => x"82f4ffc1",
  1952 => x"4cf4f6c2",
  1953 => x"6c978475",
  1954 => x"c14b494b",
  1955 => x"6a7c97a3",
  1956 => x"cc481181",
  1957 => x"66c458a6",
  1958 => x"a866c848",
  1959 => x"c087c302",
  1960 => x"66c87c97",
  1961 => x"c287c705",
  1962 => x"c448f8f6",
  1963 => x"85c178a5",
  1964 => x"04adb7c4",
  1965 => x"c487c1ff",
  1966 => x"f7c287d2",
  1967 => x"c848bfc4",
  1968 => x"cb01a8b7",
  1969 => x"02acca87",
  1970 => x"accd87c6",
  1971 => x"87f3c005",
  1972 => x"bfc4f7c2",
  1973 => x"abb7c84b",
  1974 => x"c287d203",
  1975 => x"7349c8f7",
  1976 => x"51e0c081",
  1977 => x"b7c883c1",
  1978 => x"eeff04ab",
  1979 => x"d0f7c287",
  1980 => x"50d2c148",
  1981 => x"c150cfc1",
  1982 => x"50c050cd",
  1983 => x"78c380e4",
  1984 => x"c287c9c3",
  1985 => x"49bfc4f7",
  1986 => x"c280c148",
  1987 => x"4858c8f7",
  1988 => x"7481a0c4",
  1989 => x"87f4c251",
  1990 => x"acb7f0c0",
  1991 => x"c087da04",
  1992 => x"01acb7f9",
  1993 => x"f6c287d3",
  1994 => x"ca49bffc",
  1995 => x"c04a7491",
  1996 => x"f6c28af0",
  1997 => x"a17248fc",
  1998 => x"02acca78",
  1999 => x"cd87c6c0",
  2000 => x"c7c205ac",
  2001 => x"f8f6c287",
  2002 => x"c178c348",
  2003 => x"f0c087fe",
  2004 => x"db04acb7",
  2005 => x"b7f9c087",
  2006 => x"d3c001ac",
  2007 => x"c0f7c287",
  2008 => x"91d049bf",
  2009 => x"f0c04a74",
  2010 => x"c0f7c28a",
  2011 => x"78a17248",
  2012 => x"acb7c1c1",
  2013 => x"87dbc004",
  2014 => x"acb7c6c1",
  2015 => x"87d3c001",
  2016 => x"bfc0f7c2",
  2017 => x"7491d049",
  2018 => x"8af7c04a",
  2019 => x"48c0f7c2",
  2020 => x"ca78a172",
  2021 => x"c6c002ac",
  2022 => x"05accd87",
  2023 => x"c287edc0",
  2024 => x"c348f8f6",
  2025 => x"87e4c078",
  2026 => x"05ace2c0",
  2027 => x"c087c6c0",
  2028 => x"d7c07efb",
  2029 => x"02acca87",
  2030 => x"cd87c6c0",
  2031 => x"c9c005ac",
  2032 => x"f8f6c287",
  2033 => x"c078c348",
  2034 => x"7e7487c2",
  2035 => x"d0f9026e",
  2036 => x"c3486e87",
  2037 => x"8ef499ff",
  2038 => x"4387dbf8",
  2039 => x"3d464e4f",
  2040 => x"444f4d00",
  2041 => x"4d414e00",
  2042 => x"45440045",
  2043 => x"4c554146",
  2044 => x"00303d54",
  2045 => x"00001fdb",
  2046 => x"00001fe1",
  2047 => x"00001fe5",
  2048 => x"00001fea",
  2049 => x"48d0ff1e",
  2050 => x"7178c9c8",
  2051 => x"08d4ff48",
  2052 => x"1e4f2678",
  2053 => x"eb494a71",
  2054 => x"48d0ff87",
  2055 => x"4f2678c8",
  2056 => x"711e731e",
  2057 => x"e0f7c24b",
  2058 => x"87c302bf",
  2059 => x"ff87ebc2",
  2060 => x"c9c848d0",
  2061 => x"c0497378",
  2062 => x"d4ffb1e0",
  2063 => x"c2787148",
  2064 => x"c048d4f7",
  2065 => x"0266c878",
  2066 => x"ffc387c5",
  2067 => x"c087c249",
  2068 => x"dcf7c249",
  2069 => x"0266cc59",
  2070 => x"d5c587c6",
  2071 => x"87c44ad5",
  2072 => x"4affffcf",
  2073 => x"5ae0f7c2",
  2074 => x"48e0f7c2",
  2075 => x"87c478c1",
  2076 => x"4c264d26",
  2077 => x"4f264b26",
  2078 => x"5c5b5e0e",
  2079 => x"4a710e5d",
  2080 => x"bfdcf7c2",
  2081 => x"029a724c",
  2082 => x"c84987cb",
  2083 => x"d6c0c291",
  2084 => x"c483714b",
  2085 => x"d6c4c287",
  2086 => x"134dc04b",
  2087 => x"c2997449",
  2088 => x"b9bfd8f7",
  2089 => x"7148d4ff",
  2090 => x"2cb7c178",
  2091 => x"adb7c885",
  2092 => x"c287e804",
  2093 => x"48bfd4f7",
  2094 => x"f7c280c8",
  2095 => x"effe58d8",
  2096 => x"1e731e87",
  2097 => x"4a134b71",
  2098 => x"87cb029a",
  2099 => x"e7fe4972",
  2100 => x"9a4a1387",
  2101 => x"fe87f505",
  2102 => x"c21e87da",
  2103 => x"49bfd4f7",
  2104 => x"48d4f7c2",
  2105 => x"c478a1c1",
  2106 => x"03a9b7c0",
  2107 => x"d4ff87db",
  2108 => x"d8f7c248",
  2109 => x"f7c278bf",
  2110 => x"c249bfd4",
  2111 => x"c148d4f7",
  2112 => x"c0c478a1",
  2113 => x"e504a9b7",
  2114 => x"48d0ff87",
  2115 => x"f7c278c8",
  2116 => x"78c048e0",
  2117 => x"00004f26",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"005f5f00",
  2121 => x"03000000",
  2122 => x"03030003",
  2123 => x"7f140000",
  2124 => x"7f7f147f",
  2125 => x"24000014",
  2126 => x"3a6b6b2e",
  2127 => x"6a4c0012",
  2128 => x"566c1836",
  2129 => x"7e300032",
  2130 => x"3a77594f",
  2131 => x"00004068",
  2132 => x"00030704",
  2133 => x"00000000",
  2134 => x"41633e1c",
  2135 => x"00000000",
  2136 => x"1c3e6341",
  2137 => x"2a080000",
  2138 => x"3e1c1c3e",
  2139 => x"0800082a",
  2140 => x"083e3e08",
  2141 => x"00000008",
  2142 => x"0060e080",
  2143 => x"08000000",
  2144 => x"08080808",
  2145 => x"00000008",
  2146 => x"00606000",
  2147 => x"60400000",
  2148 => x"060c1830",
  2149 => x"3e000103",
  2150 => x"7f4d597f",
  2151 => x"0400003e",
  2152 => x"007f7f06",
  2153 => x"42000000",
  2154 => x"4f597163",
  2155 => x"22000046",
  2156 => x"7f494963",
  2157 => x"1c180036",
  2158 => x"7f7f1316",
  2159 => x"27000010",
  2160 => x"7d454567",
  2161 => x"3c000039",
  2162 => x"79494b7e",
  2163 => x"01000030",
  2164 => x"0f797101",
  2165 => x"36000007",
  2166 => x"7f49497f",
  2167 => x"06000036",
  2168 => x"3f69494f",
  2169 => x"0000001e",
  2170 => x"00666600",
  2171 => x"00000000",
  2172 => x"0066e680",
  2173 => x"08000000",
  2174 => x"22141408",
  2175 => x"14000022",
  2176 => x"14141414",
  2177 => x"22000014",
  2178 => x"08141422",
  2179 => x"02000008",
  2180 => x"0f595103",
  2181 => x"7f3e0006",
  2182 => x"1f555d41",
  2183 => x"7e00001e",
  2184 => x"7f09097f",
  2185 => x"7f00007e",
  2186 => x"7f49497f",
  2187 => x"1c000036",
  2188 => x"4141633e",
  2189 => x"7f000041",
  2190 => x"3e63417f",
  2191 => x"7f00001c",
  2192 => x"4149497f",
  2193 => x"7f000041",
  2194 => x"0109097f",
  2195 => x"3e000001",
  2196 => x"7b49417f",
  2197 => x"7f00007a",
  2198 => x"7f08087f",
  2199 => x"0000007f",
  2200 => x"417f7f41",
  2201 => x"20000000",
  2202 => x"7f404060",
  2203 => x"7f7f003f",
  2204 => x"63361c08",
  2205 => x"7f000041",
  2206 => x"4040407f",
  2207 => x"7f7f0040",
  2208 => x"7f060c06",
  2209 => x"7f7f007f",
  2210 => x"7f180c06",
  2211 => x"3e00007f",
  2212 => x"7f41417f",
  2213 => x"7f00003e",
  2214 => x"0f09097f",
  2215 => x"7f3e0006",
  2216 => x"7e7f6141",
  2217 => x"7f000040",
  2218 => x"7f19097f",
  2219 => x"26000066",
  2220 => x"7b594d6f",
  2221 => x"01000032",
  2222 => x"017f7f01",
  2223 => x"3f000001",
  2224 => x"7f40407f",
  2225 => x"0f00003f",
  2226 => x"3f70703f",
  2227 => x"7f7f000f",
  2228 => x"7f301830",
  2229 => x"6341007f",
  2230 => x"361c1c36",
  2231 => x"03014163",
  2232 => x"067c7c06",
  2233 => x"71610103",
  2234 => x"43474d59",
  2235 => x"00000041",
  2236 => x"41417f7f",
  2237 => x"03010000",
  2238 => x"30180c06",
  2239 => x"00004060",
  2240 => x"7f7f4141",
  2241 => x"0c080000",
  2242 => x"0c060306",
  2243 => x"80800008",
  2244 => x"80808080",
  2245 => x"00000080",
  2246 => x"04070300",
  2247 => x"20000000",
  2248 => x"7c545474",
  2249 => x"7f000078",
  2250 => x"7c44447f",
  2251 => x"38000038",
  2252 => x"4444447c",
  2253 => x"38000000",
  2254 => x"7f44447c",
  2255 => x"3800007f",
  2256 => x"5c54547c",
  2257 => x"04000018",
  2258 => x"05057f7e",
  2259 => x"18000000",
  2260 => x"fca4a4bc",
  2261 => x"7f00007c",
  2262 => x"7c04047f",
  2263 => x"00000078",
  2264 => x"407d3d00",
  2265 => x"80000000",
  2266 => x"7dfd8080",
  2267 => x"7f000000",
  2268 => x"6c38107f",
  2269 => x"00000044",
  2270 => x"407f3f00",
  2271 => x"7c7c0000",
  2272 => x"7c0c180c",
  2273 => x"7c000078",
  2274 => x"7c04047c",
  2275 => x"38000078",
  2276 => x"7c44447c",
  2277 => x"fc000038",
  2278 => x"3c2424fc",
  2279 => x"18000018",
  2280 => x"fc24243c",
  2281 => x"7c0000fc",
  2282 => x"0c04047c",
  2283 => x"48000008",
  2284 => x"7454545c",
  2285 => x"04000020",
  2286 => x"44447f3f",
  2287 => x"3c000000",
  2288 => x"7c40407c",
  2289 => x"1c00007c",
  2290 => x"3c60603c",
  2291 => x"7c3c001c",
  2292 => x"7c603060",
  2293 => x"6c44003c",
  2294 => x"6c381038",
  2295 => x"1c000044",
  2296 => x"3c60e0bc",
  2297 => x"4400001c",
  2298 => x"4c5c7464",
  2299 => x"08000044",
  2300 => x"41773e08",
  2301 => x"00000041",
  2302 => x"007f7f00",
  2303 => x"41000000",
  2304 => x"083e7741",
  2305 => x"01020008",
  2306 => x"02020301",
  2307 => x"7f7f0001",
  2308 => x"7f7f7f7f",
  2309 => x"0808007f",
  2310 => x"3e3e1c1c",
  2311 => x"7f7f7f7f",
  2312 => x"1c1c3e3e",
  2313 => x"10000808",
  2314 => x"187c7c18",
  2315 => x"10000010",
  2316 => x"307c7c30",
  2317 => x"30100010",
  2318 => x"1e786060",
  2319 => x"66420006",
  2320 => x"663c183c",
  2321 => x"38780042",
  2322 => x"6cc6c26a",
  2323 => x"00600038",
  2324 => x"00006000",
  2325 => x"5e0e0060",
  2326 => x"0e5d5c5b",
  2327 => x"c24c711e",
  2328 => x"4dbff1f7",
  2329 => x"1ec04bc0",
  2330 => x"c702ab74",
  2331 => x"48a6c487",
  2332 => x"87c578c0",
  2333 => x"c148a6c4",
  2334 => x"1e66c478",
  2335 => x"dfee4973",
  2336 => x"c086c887",
  2337 => x"efef49e0",
  2338 => x"4aa5c487",
  2339 => x"f0f0496a",
  2340 => x"87c6f187",
  2341 => x"83c185cb",
  2342 => x"04abb7c8",
  2343 => x"2687c7ff",
  2344 => x"4c264d26",
  2345 => x"4f264b26",
  2346 => x"c24a711e",
  2347 => x"c25af5f7",
  2348 => x"c748f5f7",
  2349 => x"ddfe4978",
  2350 => x"1e4f2687",
  2351 => x"4a711e73",
  2352 => x"03aab7c0",
  2353 => x"e0c287d3",
  2354 => x"c405bfdb",
  2355 => x"c24bc187",
  2356 => x"c24bc087",
  2357 => x"c45bdfe0",
  2358 => x"dfe0c287",
  2359 => x"dbe0c25a",
  2360 => x"9ac14abf",
  2361 => x"49a2c0c1",
  2362 => x"fc87e8ec",
  2363 => x"dbe0c248",
  2364 => x"effe78bf",
  2365 => x"4a711e87",
  2366 => x"721e66c4",
  2367 => x"e9dfff49",
  2368 => x"4f262687",
  2369 => x"dbe0c21e",
  2370 => x"dcff49bf",
  2371 => x"f7c287d9",
  2372 => x"bfe848e9",
  2373 => x"e5f7c278",
  2374 => x"78bfec48",
  2375 => x"bfe9f7c2",
  2376 => x"ffc3494a",
  2377 => x"2ab7c899",
  2378 => x"b0714872",
  2379 => x"58f1f7c2",
  2380 => x"5e0e4f26",
  2381 => x"0e5d5c5b",
  2382 => x"c7ff4b71",
  2383 => x"e4f7c287",
  2384 => x"7350c048",
  2385 => x"fedbff49",
  2386 => x"4c497087",
  2387 => x"eecb9cc2",
  2388 => x"87cfcb49",
  2389 => x"c24d4970",
  2390 => x"bf97e4f7",
  2391 => x"87e4c105",
  2392 => x"c24966d0",
  2393 => x"99bfedf7",
  2394 => x"d487d705",
  2395 => x"f7c24966",
  2396 => x"0599bfe5",
  2397 => x"497387cc",
  2398 => x"87cbdbff",
  2399 => x"c1029870",
  2400 => x"4cc187c2",
  2401 => x"7587fdfd",
  2402 => x"87e3ca49",
  2403 => x"c6029870",
  2404 => x"e4f7c287",
  2405 => x"c250c148",
  2406 => x"bf97e4f7",
  2407 => x"87e4c005",
  2408 => x"bfedf7c2",
  2409 => x"9966d049",
  2410 => x"87d6ff05",
  2411 => x"bfe5f7c2",
  2412 => x"9966d449",
  2413 => x"87caff05",
  2414 => x"daff4973",
  2415 => x"987087c9",
  2416 => x"87fefe05",
  2417 => x"d7fb4874",
  2418 => x"5b5e0e87",
  2419 => x"f40e5d5c",
  2420 => x"4c4dc086",
  2421 => x"c47ebfec",
  2422 => x"f7c248a6",
  2423 => x"c178bff1",
  2424 => x"c71ec01e",
  2425 => x"87cafd49",
  2426 => x"987086c8",
  2427 => x"ff87ce02",
  2428 => x"87c7fb49",
  2429 => x"ff49dac1",
  2430 => x"c187ccd9",
  2431 => x"e4f7c24d",
  2432 => x"c302bf97",
  2433 => x"87c0c987",
  2434 => x"bfe9f7c2",
  2435 => x"dbe0c24b",
  2436 => x"ebc005bf",
  2437 => x"49fdc387",
  2438 => x"87ebd8ff",
  2439 => x"ff49fac3",
  2440 => x"7387e4d8",
  2441 => x"99ffc349",
  2442 => x"49c01e71",
  2443 => x"7387c6fb",
  2444 => x"29b7c849",
  2445 => x"49c11e71",
  2446 => x"c887fafa",
  2447 => x"87c1c686",
  2448 => x"bfedf7c2",
  2449 => x"dd029b4b",
  2450 => x"d7e0c287",
  2451 => x"dec749bf",
  2452 => x"05987087",
  2453 => x"4bc087c4",
  2454 => x"e0c287d2",
  2455 => x"87c3c749",
  2456 => x"58dbe0c2",
  2457 => x"e0c287c6",
  2458 => x"78c048d7",
  2459 => x"99c24973",
  2460 => x"c387ce05",
  2461 => x"d7ff49eb",
  2462 => x"497087cd",
  2463 => x"c20299c2",
  2464 => x"734cfb87",
  2465 => x"0599c149",
  2466 => x"f4c387ce",
  2467 => x"f6d6ff49",
  2468 => x"c2497087",
  2469 => x"87c20299",
  2470 => x"49734cfa",
  2471 => x"ce0599c8",
  2472 => x"49f5c387",
  2473 => x"87dfd6ff",
  2474 => x"99c24970",
  2475 => x"c287d502",
  2476 => x"02bff5f7",
  2477 => x"c14887ca",
  2478 => x"f9f7c288",
  2479 => x"87c2c058",
  2480 => x"4dc14cff",
  2481 => x"99c44973",
  2482 => x"c387ce05",
  2483 => x"d5ff49f2",
  2484 => x"497087f5",
  2485 => x"dc0299c2",
  2486 => x"f5f7c287",
  2487 => x"c7487ebf",
  2488 => x"c003a8b7",
  2489 => x"486e87cb",
  2490 => x"f7c280c1",
  2491 => x"c2c058f9",
  2492 => x"c14cfe87",
  2493 => x"49fdc34d",
  2494 => x"87cbd5ff",
  2495 => x"99c24970",
  2496 => x"87d5c002",
  2497 => x"bff5f7c2",
  2498 => x"87c9c002",
  2499 => x"48f5f7c2",
  2500 => x"c2c078c0",
  2501 => x"c14cfd87",
  2502 => x"49fac34d",
  2503 => x"87e7d4ff",
  2504 => x"99c24970",
  2505 => x"87d9c002",
  2506 => x"bff5f7c2",
  2507 => x"a8b7c748",
  2508 => x"87c9c003",
  2509 => x"48f5f7c2",
  2510 => x"c2c078c7",
  2511 => x"c14cfc87",
  2512 => x"acb7c04d",
  2513 => x"87d1c003",
  2514 => x"c14a66c4",
  2515 => x"026a82d8",
  2516 => x"6a87c6c0",
  2517 => x"7349744b",
  2518 => x"c31ec00f",
  2519 => x"dac11ef0",
  2520 => x"87cef749",
  2521 => x"987086c8",
  2522 => x"87e2c002",
  2523 => x"c248a6c8",
  2524 => x"78bff5f7",
  2525 => x"cb4966c8",
  2526 => x"4866c491",
  2527 => x"7e708071",
  2528 => x"c002bf6e",
  2529 => x"bf6e87c8",
  2530 => x"4966c84b",
  2531 => x"9d750f73",
  2532 => x"87c8c002",
  2533 => x"bff5f7c2",
  2534 => x"87faf249",
  2535 => x"bfdfe0c2",
  2536 => x"87ddc002",
  2537 => x"87c7c249",
  2538 => x"c0029870",
  2539 => x"f7c287d3",
  2540 => x"f249bff5",
  2541 => x"49c087e0",
  2542 => x"c287c0f4",
  2543 => x"c048dfe0",
  2544 => x"f38ef478",
  2545 => x"5e0e87da",
  2546 => x"0e5d5c5b",
  2547 => x"c24c711e",
  2548 => x"49bff1f7",
  2549 => x"4da1cdc1",
  2550 => x"6981d1c1",
  2551 => x"029c747e",
  2552 => x"a5c487cf",
  2553 => x"c27b744b",
  2554 => x"49bff1f7",
  2555 => x"6e87f9f2",
  2556 => x"059c747b",
  2557 => x"4bc087c4",
  2558 => x"4bc187c2",
  2559 => x"faf24973",
  2560 => x"0266d487",
  2561 => x"da4987c7",
  2562 => x"c24a7087",
  2563 => x"c24ac087",
  2564 => x"265ae3e0",
  2565 => x"0087c9f2",
  2566 => x"00000000",
  2567 => x"00000000",
  2568 => x"1e000000",
  2569 => x"c8ff4a71",
  2570 => x"a17249bf",
  2571 => x"1e4f2648",
  2572 => x"89bfc8ff",
  2573 => x"c0c0c0fe",
  2574 => x"01a9c0c0",
  2575 => x"4ac087c4",
  2576 => x"4ac187c2",
  2577 => x"4f264872",
  2578 => x"d6e2c21e",
  2579 => x"b9c149bf",
  2580 => x"59dae2c2",
  2581 => x"c348d4ff",
  2582 => x"d0ff78ff",
  2583 => x"78e1c048",
  2584 => x"c148d4ff",
  2585 => x"7131c478",
  2586 => x"48d0ff78",
  2587 => x"2678e0c0",
  2588 => x"e2c21e4f",
  2589 => x"f2c21eca",
  2590 => x"fcfd49d8",
  2591 => x"86c487c7",
  2592 => x"c3029870",
  2593 => x"87c0ff87",
  2594 => x"35314f26",
  2595 => x"205a484b",
  2596 => x"46432020",
  2597 => x"00000047",
  2598 => x"5e0e0000",
  2599 => x"0e5d5c5b",
  2600 => x"bfe5f7c2",
  2601 => x"c3e4c24a",
  2602 => x"724c49bf",
  2603 => x"ff4d71bc",
  2604 => x"c087ebc6",
  2605 => x"d049744b",
  2606 => x"e7c00299",
  2607 => x"48d0ff87",
  2608 => x"ff78e1c8",
  2609 => x"78c548d4",
  2610 => x"99d04975",
  2611 => x"c387c302",
  2612 => x"e4c278f0",
  2613 => x"817349f1",
  2614 => x"d4ff4811",
  2615 => x"d0ff7808",
  2616 => x"78e0c048",
  2617 => x"832d2cc1",
  2618 => x"ff04abc8",
  2619 => x"c5ff87c7",
  2620 => x"e4c287e4",
  2621 => x"f7c248c3",
  2622 => x"2678bfe5",
  2623 => x"264c264d",
  2624 => x"004f264b",
  2625 => x"1e000000",
  2626 => x"48c9e7c1",
  2627 => x"e4c250de",
  2628 => x"d9fe49da",
  2629 => x"48c087f1",
  2630 => x"544a4f26",
  2631 => x"5254554f",
  2632 => x"52414e55",
  2633 => x"f21e0043",
  2634 => x"edfd87df",
  2635 => x"2687f887",
  2636 => x"261e164f",
  2637 => x"3d362e25",
  2638 => x"3d362e3e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
