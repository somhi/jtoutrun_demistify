
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d8",x"fa",x"c2",x"87"),
    12 => (x"86",x"c0",x"c5",x"4e"),
    13 => (x"49",x"d8",x"fa",x"c2"),
    14 => (x"48",x"cc",x"e7",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"f4",x"e5"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"71",x"1e",x"4f",x"26"),
    53 => (x"49",x"66",x"c4",x"4a"),
    54 => (x"c8",x"88",x"c1",x"48"),
    55 => (x"99",x"71",x"58",x"a6"),
    56 => (x"ff",x"87",x"d6",x"02"),
    57 => (x"ff",x"c3",x"48",x"d4"),
    58 => (x"c4",x"52",x"68",x"78"),
    59 => (x"c1",x"48",x"49",x"66"),
    60 => (x"58",x"a6",x"c8",x"88"),
    61 => (x"ea",x"05",x"99",x"71"),
    62 => (x"1e",x"4f",x"26",x"87"),
    63 => (x"d4",x"ff",x"1e",x"73"),
    64 => (x"7b",x"ff",x"c3",x"4b"),
    65 => (x"ff",x"c3",x"4a",x"6b"),
    66 => (x"c8",x"49",x"6b",x"7b"),
    67 => (x"c3",x"b1",x"72",x"32"),
    68 => (x"4a",x"6b",x"7b",x"ff"),
    69 => (x"b2",x"71",x"31",x"c8"),
    70 => (x"6b",x"7b",x"ff",x"c3"),
    71 => (x"72",x"32",x"c8",x"49"),
    72 => (x"c4",x"48",x"71",x"b1"),
    73 => (x"26",x"4d",x"26",x"87"),
    74 => (x"26",x"4b",x"26",x"4c"),
    75 => (x"5b",x"5e",x"0e",x"4f"),
    76 => (x"71",x"0e",x"5d",x"5c"),
    77 => (x"4c",x"d4",x"ff",x"4a"),
    78 => (x"ff",x"c3",x"49",x"72"),
    79 => (x"c2",x"7c",x"71",x"99"),
    80 => (x"05",x"bf",x"cc",x"e7"),
    81 => (x"66",x"d0",x"87",x"c8"),
    82 => (x"d4",x"30",x"c9",x"48"),
    83 => (x"66",x"d0",x"58",x"a6"),
    84 => (x"c3",x"29",x"d8",x"49"),
    85 => (x"7c",x"71",x"99",x"ff"),
    86 => (x"d0",x"49",x"66",x"d0"),
    87 => (x"99",x"ff",x"c3",x"29"),
    88 => (x"66",x"d0",x"7c",x"71"),
    89 => (x"c3",x"29",x"c8",x"49"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"c3",x"49",x"66",x"d0"),
    92 => (x"7c",x"71",x"99",x"ff"),
    93 => (x"29",x"d0",x"49",x"72"),
    94 => (x"71",x"99",x"ff",x"c3"),
    95 => (x"c9",x"4b",x"6c",x"7c"),
    96 => (x"c3",x"4d",x"ff",x"f0"),
    97 => (x"d0",x"05",x"ab",x"ff"),
    98 => (x"7c",x"ff",x"c3",x"87"),
    99 => (x"8d",x"c1",x"4b",x"6c"),
   100 => (x"c3",x"87",x"c6",x"02"),
   101 => (x"f0",x"02",x"ab",x"ff"),
   102 => (x"fe",x"48",x"73",x"87"),
   103 => (x"c0",x"1e",x"87",x"c7"),
   104 => (x"48",x"d4",x"ff",x"49"),
   105 => (x"c1",x"78",x"ff",x"c3"),
   106 => (x"b7",x"c8",x"c3",x"81"),
   107 => (x"87",x"f1",x"04",x"a9"),
   108 => (x"73",x"1e",x"4f",x"26"),
   109 => (x"c4",x"87",x"e7",x"1e"),
   110 => (x"c0",x"4b",x"df",x"f8"),
   111 => (x"f0",x"ff",x"c0",x"1e"),
   112 => (x"fd",x"49",x"f7",x"c1"),
   113 => (x"86",x"c4",x"87",x"e7"),
   114 => (x"c0",x"05",x"a8",x"c1"),
   115 => (x"d4",x"ff",x"87",x"ea"),
   116 => (x"78",x"ff",x"c3",x"48"),
   117 => (x"c0",x"c0",x"c0",x"c1"),
   118 => (x"c0",x"1e",x"c0",x"c0"),
   119 => (x"e9",x"c1",x"f0",x"e1"),
   120 => (x"87",x"c9",x"fd",x"49"),
   121 => (x"98",x"70",x"86",x"c4"),
   122 => (x"ff",x"87",x"ca",x"05"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"cb",x"48",x"c1",x"78"),
   125 => (x"87",x"e6",x"fe",x"87"),
   126 => (x"fe",x"05",x"8b",x"c1"),
   127 => (x"48",x"c0",x"87",x"fd"),
   128 => (x"1e",x"87",x"e6",x"fc"),
   129 => (x"d4",x"ff",x"1e",x"73"),
   130 => (x"78",x"ff",x"c3",x"48"),
   131 => (x"1e",x"c0",x"4b",x"d3"),
   132 => (x"c1",x"f0",x"ff",x"c0"),
   133 => (x"d4",x"fc",x"49",x"c1"),
   134 => (x"70",x"86",x"c4",x"87"),
   135 => (x"87",x"ca",x"05",x"98"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"48",x"c1",x"78",x"ff"),
   138 => (x"f1",x"fd",x"87",x"cb"),
   139 => (x"05",x"8b",x"c1",x"87"),
   140 => (x"c0",x"87",x"db",x"ff"),
   141 => (x"87",x"f1",x"fb",x"48"),
   142 => (x"5c",x"5b",x"5e",x"0e"),
   143 => (x"4c",x"d4",x"ff",x"0e"),
   144 => (x"c6",x"87",x"db",x"fd"),
   145 => (x"e1",x"c0",x"1e",x"ea"),
   146 => (x"49",x"c8",x"c1",x"f0"),
   147 => (x"c4",x"87",x"de",x"fb"),
   148 => (x"02",x"a8",x"c1",x"86"),
   149 => (x"ea",x"fe",x"87",x"c8"),
   150 => (x"c1",x"48",x"c0",x"87"),
   151 => (x"da",x"fa",x"87",x"e2"),
   152 => (x"cf",x"49",x"70",x"87"),
   153 => (x"c6",x"99",x"ff",x"ff"),
   154 => (x"c8",x"02",x"a9",x"ea"),
   155 => (x"87",x"d3",x"fe",x"87"),
   156 => (x"cb",x"c1",x"48",x"c0"),
   157 => (x"7c",x"ff",x"c3",x"87"),
   158 => (x"fc",x"4b",x"f1",x"c0"),
   159 => (x"98",x"70",x"87",x"f4"),
   160 => (x"87",x"eb",x"c0",x"02"),
   161 => (x"ff",x"c0",x"1e",x"c0"),
   162 => (x"49",x"fa",x"c1",x"f0"),
   163 => (x"c4",x"87",x"de",x"fa"),
   164 => (x"05",x"98",x"70",x"86"),
   165 => (x"ff",x"c3",x"87",x"d9"),
   166 => (x"c3",x"49",x"6c",x"7c"),
   167 => (x"7c",x"7c",x"7c",x"ff"),
   168 => (x"99",x"c0",x"c1",x"7c"),
   169 => (x"c1",x"87",x"c4",x"02"),
   170 => (x"c0",x"87",x"d5",x"48"),
   171 => (x"c2",x"87",x"d1",x"48"),
   172 => (x"87",x"c4",x"05",x"ab"),
   173 => (x"87",x"c8",x"48",x"c0"),
   174 => (x"fe",x"05",x"8b",x"c1"),
   175 => (x"48",x"c0",x"87",x"fd"),
   176 => (x"1e",x"87",x"e4",x"f9"),
   177 => (x"e7",x"c2",x"1e",x"73"),
   178 => (x"78",x"c1",x"48",x"cc"),
   179 => (x"d0",x"ff",x"4b",x"c7"),
   180 => (x"fb",x"78",x"c2",x"48"),
   181 => (x"d0",x"ff",x"87",x"c8"),
   182 => (x"c0",x"78",x"c3",x"48"),
   183 => (x"d0",x"e5",x"c0",x"1e"),
   184 => (x"f9",x"49",x"c0",x"c1"),
   185 => (x"86",x"c4",x"87",x"c7"),
   186 => (x"c1",x"05",x"a8",x"c1"),
   187 => (x"ab",x"c2",x"4b",x"87"),
   188 => (x"c0",x"87",x"c5",x"05"),
   189 => (x"87",x"f9",x"c0",x"48"),
   190 => (x"ff",x"05",x"8b",x"c1"),
   191 => (x"f7",x"fc",x"87",x"d0"),
   192 => (x"d0",x"e7",x"c2",x"87"),
   193 => (x"05",x"98",x"70",x"58"),
   194 => (x"1e",x"c1",x"87",x"cd"),
   195 => (x"c1",x"f0",x"ff",x"c0"),
   196 => (x"d8",x"f8",x"49",x"d0"),
   197 => (x"ff",x"86",x"c4",x"87"),
   198 => (x"ff",x"c3",x"48",x"d4"),
   199 => (x"87",x"fc",x"c2",x"78"),
   200 => (x"58",x"d4",x"e7",x"c2"),
   201 => (x"c2",x"48",x"d0",x"ff"),
   202 => (x"48",x"d4",x"ff",x"78"),
   203 => (x"c1",x"78",x"ff",x"c3"),
   204 => (x"87",x"f5",x"f7",x"48"),
   205 => (x"5c",x"5b",x"5e",x"0e"),
   206 => (x"4b",x"71",x"0e",x"5d"),
   207 => (x"ee",x"c5",x"4c",x"c0"),
   208 => (x"ff",x"4a",x"df",x"cd"),
   209 => (x"ff",x"c3",x"48",x"d4"),
   210 => (x"c3",x"49",x"68",x"78"),
   211 => (x"c0",x"05",x"a9",x"fe"),
   212 => (x"4d",x"70",x"87",x"fd"),
   213 => (x"cc",x"02",x"9b",x"73"),
   214 => (x"1e",x"66",x"d0",x"87"),
   215 => (x"f1",x"f5",x"49",x"73"),
   216 => (x"d6",x"86",x"c4",x"87"),
   217 => (x"48",x"d0",x"ff",x"87"),
   218 => (x"c3",x"78",x"d1",x"c4"),
   219 => (x"66",x"d0",x"7d",x"ff"),
   220 => (x"d4",x"88",x"c1",x"48"),
   221 => (x"98",x"70",x"58",x"a6"),
   222 => (x"ff",x"87",x"f0",x"05"),
   223 => (x"ff",x"c3",x"48",x"d4"),
   224 => (x"9b",x"73",x"78",x"78"),
   225 => (x"ff",x"87",x"c5",x"05"),
   226 => (x"78",x"d0",x"48",x"d0"),
   227 => (x"c1",x"4c",x"4a",x"c1"),
   228 => (x"ee",x"fe",x"05",x"8a"),
   229 => (x"f6",x"48",x"74",x"87"),
   230 => (x"73",x"1e",x"87",x"cb"),
   231 => (x"c0",x"4a",x"71",x"1e"),
   232 => (x"48",x"d4",x"ff",x"4b"),
   233 => (x"ff",x"78",x"ff",x"c3"),
   234 => (x"c3",x"c4",x"48",x"d0"),
   235 => (x"48",x"d4",x"ff",x"78"),
   236 => (x"72",x"78",x"ff",x"c3"),
   237 => (x"f0",x"ff",x"c0",x"1e"),
   238 => (x"f5",x"49",x"d1",x"c1"),
   239 => (x"86",x"c4",x"87",x"ef"),
   240 => (x"d2",x"05",x"98",x"70"),
   241 => (x"1e",x"c0",x"c8",x"87"),
   242 => (x"fd",x"49",x"66",x"cc"),
   243 => (x"86",x"c4",x"87",x"e6"),
   244 => (x"d0",x"ff",x"4b",x"70"),
   245 => (x"73",x"78",x"c2",x"48"),
   246 => (x"87",x"cd",x"f5",x"48"),
   247 => (x"5c",x"5b",x"5e",x"0e"),
   248 => (x"1e",x"c0",x"0e",x"5d"),
   249 => (x"c1",x"f0",x"ff",x"c0"),
   250 => (x"c0",x"f5",x"49",x"c9"),
   251 => (x"c2",x"1e",x"d2",x"87"),
   252 => (x"fc",x"49",x"d4",x"e7"),
   253 => (x"86",x"c8",x"87",x"fe"),
   254 => (x"84",x"c1",x"4c",x"c0"),
   255 => (x"04",x"ac",x"b7",x"d2"),
   256 => (x"e7",x"c2",x"87",x"f8"),
   257 => (x"49",x"bf",x"97",x"d4"),
   258 => (x"c1",x"99",x"c0",x"c3"),
   259 => (x"c0",x"05",x"a9",x"c0"),
   260 => (x"e7",x"c2",x"87",x"e7"),
   261 => (x"49",x"bf",x"97",x"db"),
   262 => (x"e7",x"c2",x"31",x"d0"),
   263 => (x"4a",x"bf",x"97",x"dc"),
   264 => (x"b1",x"72",x"32",x"c8"),
   265 => (x"97",x"dd",x"e7",x"c2"),
   266 => (x"71",x"b1",x"4a",x"bf"),
   267 => (x"ff",x"ff",x"cf",x"4c"),
   268 => (x"84",x"c1",x"9c",x"ff"),
   269 => (x"e7",x"c1",x"34",x"ca"),
   270 => (x"dd",x"e7",x"c2",x"87"),
   271 => (x"c1",x"49",x"bf",x"97"),
   272 => (x"c2",x"99",x"c6",x"31"),
   273 => (x"bf",x"97",x"de",x"e7"),
   274 => (x"2a",x"b7",x"c7",x"4a"),
   275 => (x"e7",x"c2",x"b1",x"72"),
   276 => (x"4a",x"bf",x"97",x"d9"),
   277 => (x"c2",x"9d",x"cf",x"4d"),
   278 => (x"bf",x"97",x"da",x"e7"),
   279 => (x"ca",x"9a",x"c3",x"4a"),
   280 => (x"db",x"e7",x"c2",x"32"),
   281 => (x"c2",x"4b",x"bf",x"97"),
   282 => (x"c2",x"b2",x"73",x"33"),
   283 => (x"bf",x"97",x"dc",x"e7"),
   284 => (x"9b",x"c0",x"c3",x"4b"),
   285 => (x"73",x"2b",x"b7",x"c6"),
   286 => (x"c1",x"81",x"c2",x"b2"),
   287 => (x"70",x"30",x"71",x"48"),
   288 => (x"75",x"48",x"c1",x"49"),
   289 => (x"72",x"4d",x"70",x"30"),
   290 => (x"71",x"84",x"c1",x"4c"),
   291 => (x"b7",x"c0",x"c8",x"94"),
   292 => (x"87",x"cc",x"06",x"ad"),
   293 => (x"2d",x"b7",x"34",x"c1"),
   294 => (x"ad",x"b7",x"c0",x"c8"),
   295 => (x"87",x"f4",x"ff",x"01"),
   296 => (x"c0",x"f2",x"48",x"74"),
   297 => (x"5b",x"5e",x"0e",x"87"),
   298 => (x"f8",x"0e",x"5d",x"5c"),
   299 => (x"fa",x"ef",x"c2",x"86"),
   300 => (x"c2",x"78",x"c0",x"48"),
   301 => (x"c0",x"1e",x"f2",x"e7"),
   302 => (x"87",x"de",x"fb",x"49"),
   303 => (x"98",x"70",x"86",x"c4"),
   304 => (x"c0",x"87",x"c5",x"05"),
   305 => (x"87",x"ce",x"c9",x"48"),
   306 => (x"7e",x"c1",x"4d",x"c0"),
   307 => (x"bf",x"e2",x"f5",x"c0"),
   308 => (x"e8",x"e8",x"c2",x"49"),
   309 => (x"4b",x"c8",x"71",x"4a"),
   310 => (x"70",x"87",x"cf",x"ee"),
   311 => (x"87",x"c2",x"05",x"98"),
   312 => (x"f5",x"c0",x"7e",x"c0"),
   313 => (x"c2",x"49",x"bf",x"de"),
   314 => (x"71",x"4a",x"c4",x"e9"),
   315 => (x"f9",x"ed",x"4b",x"c8"),
   316 => (x"05",x"98",x"70",x"87"),
   317 => (x"7e",x"c0",x"87",x"c2"),
   318 => (x"fd",x"c0",x"02",x"6e"),
   319 => (x"f8",x"ee",x"c2",x"87"),
   320 => (x"ef",x"c2",x"4d",x"bf"),
   321 => (x"7e",x"bf",x"9f",x"f0"),
   322 => (x"ea",x"d6",x"c5",x"48"),
   323 => (x"87",x"c7",x"05",x"a8"),
   324 => (x"bf",x"f8",x"ee",x"c2"),
   325 => (x"6e",x"87",x"ce",x"4d"),
   326 => (x"d5",x"e9",x"ca",x"48"),
   327 => (x"87",x"c5",x"02",x"a8"),
   328 => (x"f1",x"c7",x"48",x"c0"),
   329 => (x"f2",x"e7",x"c2",x"87"),
   330 => (x"f9",x"49",x"75",x"1e"),
   331 => (x"86",x"c4",x"87",x"ec"),
   332 => (x"c5",x"05",x"98",x"70"),
   333 => (x"c7",x"48",x"c0",x"87"),
   334 => (x"f5",x"c0",x"87",x"dc"),
   335 => (x"c2",x"49",x"bf",x"de"),
   336 => (x"71",x"4a",x"c4",x"e9"),
   337 => (x"e1",x"ec",x"4b",x"c8"),
   338 => (x"05",x"98",x"70",x"87"),
   339 => (x"ef",x"c2",x"87",x"c8"),
   340 => (x"78",x"c1",x"48",x"fa"),
   341 => (x"f5",x"c0",x"87",x"da"),
   342 => (x"c2",x"49",x"bf",x"e2"),
   343 => (x"71",x"4a",x"e8",x"e8"),
   344 => (x"c5",x"ec",x"4b",x"c8"),
   345 => (x"02",x"98",x"70",x"87"),
   346 => (x"c0",x"87",x"c5",x"c0"),
   347 => (x"87",x"e6",x"c6",x"48"),
   348 => (x"97",x"f0",x"ef",x"c2"),
   349 => (x"d5",x"c1",x"49",x"bf"),
   350 => (x"cd",x"c0",x"05",x"a9"),
   351 => (x"f1",x"ef",x"c2",x"87"),
   352 => (x"c2",x"49",x"bf",x"97"),
   353 => (x"c0",x"02",x"a9",x"ea"),
   354 => (x"48",x"c0",x"87",x"c5"),
   355 => (x"c2",x"87",x"c7",x"c6"),
   356 => (x"bf",x"97",x"f2",x"e7"),
   357 => (x"e9",x"c3",x"48",x"7e"),
   358 => (x"ce",x"c0",x"02",x"a8"),
   359 => (x"c3",x"48",x"6e",x"87"),
   360 => (x"c0",x"02",x"a8",x"eb"),
   361 => (x"48",x"c0",x"87",x"c5"),
   362 => (x"c2",x"87",x"eb",x"c5"),
   363 => (x"bf",x"97",x"fd",x"e7"),
   364 => (x"c0",x"05",x"99",x"49"),
   365 => (x"e7",x"c2",x"87",x"cc"),
   366 => (x"49",x"bf",x"97",x"fe"),
   367 => (x"c0",x"02",x"a9",x"c2"),
   368 => (x"48",x"c0",x"87",x"c5"),
   369 => (x"c2",x"87",x"cf",x"c5"),
   370 => (x"bf",x"97",x"ff",x"e7"),
   371 => (x"f6",x"ef",x"c2",x"48"),
   372 => (x"48",x"4c",x"70",x"58"),
   373 => (x"ef",x"c2",x"88",x"c1"),
   374 => (x"e8",x"c2",x"58",x"fa"),
   375 => (x"49",x"bf",x"97",x"c0"),
   376 => (x"e8",x"c2",x"81",x"75"),
   377 => (x"4a",x"bf",x"97",x"c1"),
   378 => (x"a1",x"72",x"32",x"c8"),
   379 => (x"c7",x"f4",x"c2",x"7e"),
   380 => (x"c2",x"78",x"6e",x"48"),
   381 => (x"bf",x"97",x"c2",x"e8"),
   382 => (x"58",x"a6",x"c8",x"48"),
   383 => (x"bf",x"fa",x"ef",x"c2"),
   384 => (x"87",x"d4",x"c2",x"02"),
   385 => (x"bf",x"de",x"f5",x"c0"),
   386 => (x"c4",x"e9",x"c2",x"49"),
   387 => (x"4b",x"c8",x"71",x"4a"),
   388 => (x"70",x"87",x"d7",x"e9"),
   389 => (x"c5",x"c0",x"02",x"98"),
   390 => (x"c3",x"48",x"c0",x"87"),
   391 => (x"ef",x"c2",x"87",x"f8"),
   392 => (x"c2",x"4c",x"bf",x"f2"),
   393 => (x"c2",x"5c",x"db",x"f4"),
   394 => (x"bf",x"97",x"d7",x"e8"),
   395 => (x"c2",x"31",x"c8",x"49"),
   396 => (x"bf",x"97",x"d6",x"e8"),
   397 => (x"c2",x"49",x"a1",x"4a"),
   398 => (x"bf",x"97",x"d8",x"e8"),
   399 => (x"72",x"32",x"d0",x"4a"),
   400 => (x"e8",x"c2",x"49",x"a1"),
   401 => (x"4a",x"bf",x"97",x"d9"),
   402 => (x"a1",x"72",x"32",x"d8"),
   403 => (x"91",x"66",x"c4",x"49"),
   404 => (x"bf",x"c7",x"f4",x"c2"),
   405 => (x"cf",x"f4",x"c2",x"81"),
   406 => (x"df",x"e8",x"c2",x"59"),
   407 => (x"c8",x"4a",x"bf",x"97"),
   408 => (x"de",x"e8",x"c2",x"32"),
   409 => (x"a2",x"4b",x"bf",x"97"),
   410 => (x"e0",x"e8",x"c2",x"4a"),
   411 => (x"d0",x"4b",x"bf",x"97"),
   412 => (x"4a",x"a2",x"73",x"33"),
   413 => (x"97",x"e1",x"e8",x"c2"),
   414 => (x"9b",x"cf",x"4b",x"bf"),
   415 => (x"a2",x"73",x"33",x"d8"),
   416 => (x"d3",x"f4",x"c2",x"4a"),
   417 => (x"cf",x"f4",x"c2",x"5a"),
   418 => (x"8a",x"c2",x"4a",x"bf"),
   419 => (x"f4",x"c2",x"92",x"74"),
   420 => (x"a1",x"72",x"48",x"d3"),
   421 => (x"87",x"ca",x"c1",x"78"),
   422 => (x"97",x"c4",x"e8",x"c2"),
   423 => (x"31",x"c8",x"49",x"bf"),
   424 => (x"97",x"c3",x"e8",x"c2"),
   425 => (x"49",x"a1",x"4a",x"bf"),
   426 => (x"59",x"c2",x"f0",x"c2"),
   427 => (x"bf",x"fe",x"ef",x"c2"),
   428 => (x"c7",x"31",x"c5",x"49"),
   429 => (x"29",x"c9",x"81",x"ff"),
   430 => (x"59",x"db",x"f4",x"c2"),
   431 => (x"97",x"c9",x"e8",x"c2"),
   432 => (x"32",x"c8",x"4a",x"bf"),
   433 => (x"97",x"c8",x"e8",x"c2"),
   434 => (x"4a",x"a2",x"4b",x"bf"),
   435 => (x"6e",x"92",x"66",x"c4"),
   436 => (x"d7",x"f4",x"c2",x"82"),
   437 => (x"cf",x"f4",x"c2",x"5a"),
   438 => (x"c2",x"78",x"c0",x"48"),
   439 => (x"72",x"48",x"cb",x"f4"),
   440 => (x"f4",x"c2",x"78",x"a1"),
   441 => (x"f4",x"c2",x"48",x"db"),
   442 => (x"c2",x"78",x"bf",x"cf"),
   443 => (x"c2",x"48",x"df",x"f4"),
   444 => (x"78",x"bf",x"d3",x"f4"),
   445 => (x"bf",x"fa",x"ef",x"c2"),
   446 => (x"87",x"c9",x"c0",x"02"),
   447 => (x"30",x"c4",x"48",x"74"),
   448 => (x"c9",x"c0",x"7e",x"70"),
   449 => (x"d7",x"f4",x"c2",x"87"),
   450 => (x"30",x"c4",x"48",x"bf"),
   451 => (x"ef",x"c2",x"7e",x"70"),
   452 => (x"78",x"6e",x"48",x"fe"),
   453 => (x"8e",x"f8",x"48",x"c1"),
   454 => (x"4c",x"26",x"4d",x"26"),
   455 => (x"4f",x"26",x"4b",x"26"),
   456 => (x"5c",x"5b",x"5e",x"0e"),
   457 => (x"4a",x"71",x"0e",x"5d"),
   458 => (x"bf",x"fa",x"ef",x"c2"),
   459 => (x"72",x"87",x"cb",x"02"),
   460 => (x"72",x"2b",x"c7",x"4b"),
   461 => (x"9c",x"ff",x"c1",x"4c"),
   462 => (x"4b",x"72",x"87",x"c9"),
   463 => (x"4c",x"72",x"2b",x"c8"),
   464 => (x"c2",x"9c",x"ff",x"c3"),
   465 => (x"83",x"bf",x"c7",x"f4"),
   466 => (x"bf",x"da",x"f5",x"c0"),
   467 => (x"87",x"d9",x"02",x"ab"),
   468 => (x"5b",x"de",x"f5",x"c0"),
   469 => (x"1e",x"f2",x"e7",x"c2"),
   470 => (x"fd",x"f0",x"49",x"73"),
   471 => (x"70",x"86",x"c4",x"87"),
   472 => (x"87",x"c5",x"05",x"98"),
   473 => (x"e6",x"c0",x"48",x"c0"),
   474 => (x"fa",x"ef",x"c2",x"87"),
   475 => (x"87",x"d2",x"02",x"bf"),
   476 => (x"91",x"c4",x"49",x"74"),
   477 => (x"81",x"f2",x"e7",x"c2"),
   478 => (x"ff",x"cf",x"4d",x"69"),
   479 => (x"9d",x"ff",x"ff",x"ff"),
   480 => (x"49",x"74",x"87",x"cb"),
   481 => (x"e7",x"c2",x"91",x"c2"),
   482 => (x"69",x"9f",x"81",x"f2"),
   483 => (x"fe",x"48",x"75",x"4d"),
   484 => (x"5e",x"0e",x"87",x"c6"),
   485 => (x"0e",x"5d",x"5c",x"5b"),
   486 => (x"c0",x"4d",x"71",x"1e"),
   487 => (x"cf",x"49",x"c1",x"1e"),
   488 => (x"86",x"c4",x"87",x"dc"),
   489 => (x"02",x"9c",x"4c",x"70"),
   490 => (x"c2",x"87",x"c0",x"c1"),
   491 => (x"75",x"4a",x"c2",x"f0"),
   492 => (x"87",x"db",x"e2",x"49"),
   493 => (x"c0",x"02",x"98",x"70"),
   494 => (x"4a",x"74",x"87",x"f1"),
   495 => (x"4b",x"cb",x"49",x"75"),
   496 => (x"70",x"87",x"c1",x"e3"),
   497 => (x"e2",x"c0",x"02",x"98"),
   498 => (x"74",x"1e",x"c0",x"87"),
   499 => (x"87",x"c7",x"02",x"9c"),
   500 => (x"c0",x"48",x"a6",x"c4"),
   501 => (x"c4",x"87",x"c5",x"78"),
   502 => (x"78",x"c1",x"48",x"a6"),
   503 => (x"ce",x"49",x"66",x"c4"),
   504 => (x"86",x"c4",x"87",x"dc"),
   505 => (x"05",x"9c",x"4c",x"70"),
   506 => (x"74",x"87",x"c0",x"ff"),
   507 => (x"e7",x"fc",x"26",x"48"),
   508 => (x"5b",x"5e",x"0e",x"87"),
   509 => (x"1e",x"0e",x"5d",x"5c"),
   510 => (x"05",x"9b",x"4b",x"71"),
   511 => (x"48",x"c0",x"87",x"c5"),
   512 => (x"c8",x"87",x"e5",x"c1"),
   513 => (x"7d",x"c0",x"4d",x"a3"),
   514 => (x"c7",x"02",x"66",x"d4"),
   515 => (x"97",x"66",x"d4",x"87"),
   516 => (x"87",x"c5",x"05",x"bf"),
   517 => (x"cf",x"c1",x"48",x"c0"),
   518 => (x"49",x"66",x"d4",x"87"),
   519 => (x"70",x"87",x"f3",x"fd"),
   520 => (x"c1",x"02",x"9c",x"4c"),
   521 => (x"a4",x"dc",x"87",x"c0"),
   522 => (x"da",x"7d",x"69",x"49"),
   523 => (x"a3",x"c4",x"49",x"a4"),
   524 => (x"7a",x"69",x"9f",x"4a"),
   525 => (x"bf",x"fa",x"ef",x"c2"),
   526 => (x"d4",x"87",x"d2",x"02"),
   527 => (x"69",x"9f",x"49",x"a4"),
   528 => (x"ff",x"ff",x"c0",x"49"),
   529 => (x"d0",x"48",x"71",x"99"),
   530 => (x"c2",x"7e",x"70",x"30"),
   531 => (x"6e",x"7e",x"c0",x"87"),
   532 => (x"80",x"6a",x"48",x"49"),
   533 => (x"7b",x"c0",x"7a",x"70"),
   534 => (x"6a",x"49",x"a3",x"cc"),
   535 => (x"49",x"a3",x"d0",x"79"),
   536 => (x"48",x"c1",x"79",x"c0"),
   537 => (x"48",x"c0",x"87",x"c2"),
   538 => (x"87",x"ec",x"fa",x"26"),
   539 => (x"5c",x"5b",x"5e",x"0e"),
   540 => (x"4c",x"71",x"0e",x"5d"),
   541 => (x"ca",x"c1",x"02",x"9c"),
   542 => (x"49",x"a4",x"c8",x"87"),
   543 => (x"c2",x"c1",x"02",x"69"),
   544 => (x"4a",x"66",x"d0",x"87"),
   545 => (x"d4",x"82",x"49",x"6c"),
   546 => (x"66",x"d0",x"5a",x"a6"),
   547 => (x"ef",x"c2",x"b9",x"4d"),
   548 => (x"ff",x"4a",x"bf",x"f6"),
   549 => (x"71",x"99",x"72",x"ba"),
   550 => (x"e4",x"c0",x"02",x"99"),
   551 => (x"4b",x"a4",x"c4",x"87"),
   552 => (x"fb",x"f9",x"49",x"6b"),
   553 => (x"c2",x"7b",x"70",x"87"),
   554 => (x"49",x"bf",x"f2",x"ef"),
   555 => (x"7c",x"71",x"81",x"6c"),
   556 => (x"ef",x"c2",x"b9",x"75"),
   557 => (x"ff",x"4a",x"bf",x"f6"),
   558 => (x"71",x"99",x"72",x"ba"),
   559 => (x"dc",x"ff",x"05",x"99"),
   560 => (x"f9",x"7c",x"75",x"87"),
   561 => (x"73",x"1e",x"87",x"d2"),
   562 => (x"9b",x"4b",x"71",x"1e"),
   563 => (x"c8",x"87",x"c7",x"02"),
   564 => (x"05",x"69",x"49",x"a3"),
   565 => (x"48",x"c0",x"87",x"c5"),
   566 => (x"c2",x"87",x"f7",x"c0"),
   567 => (x"4a",x"bf",x"cb",x"f4"),
   568 => (x"69",x"49",x"a3",x"c4"),
   569 => (x"c2",x"89",x"c2",x"49"),
   570 => (x"91",x"bf",x"f2",x"ef"),
   571 => (x"c2",x"4a",x"a2",x"71"),
   572 => (x"49",x"bf",x"f6",x"ef"),
   573 => (x"a2",x"71",x"99",x"6b"),
   574 => (x"de",x"f5",x"c0",x"4a"),
   575 => (x"1e",x"66",x"c8",x"5a"),
   576 => (x"d5",x"ea",x"49",x"72"),
   577 => (x"70",x"86",x"c4",x"87"),
   578 => (x"87",x"c4",x"05",x"98"),
   579 => (x"87",x"c2",x"48",x"c0"),
   580 => (x"c7",x"f8",x"48",x"c1"),
   581 => (x"5b",x"5e",x"0e",x"87"),
   582 => (x"1e",x"0e",x"5d",x"5c"),
   583 => (x"66",x"d4",x"4b",x"71"),
   584 => (x"73",x"2c",x"c9",x"4c"),
   585 => (x"cf",x"c1",x"02",x"9b"),
   586 => (x"49",x"a3",x"c8",x"87"),
   587 => (x"c7",x"c1",x"02",x"69"),
   588 => (x"4d",x"a3",x"d0",x"87"),
   589 => (x"c2",x"7d",x"66",x"d4"),
   590 => (x"49",x"bf",x"f6",x"ef"),
   591 => (x"4a",x"6b",x"b9",x"ff"),
   592 => (x"ac",x"71",x"7e",x"99"),
   593 => (x"c0",x"87",x"cd",x"03"),
   594 => (x"a3",x"cc",x"7d",x"7b"),
   595 => (x"49",x"a3",x"c4",x"4a"),
   596 => (x"87",x"c2",x"79",x"6a"),
   597 => (x"9c",x"74",x"8c",x"72"),
   598 => (x"49",x"87",x"dd",x"02"),
   599 => (x"fc",x"49",x"73",x"1e"),
   600 => (x"86",x"c4",x"87",x"ca"),
   601 => (x"c7",x"49",x"66",x"d4"),
   602 => (x"cb",x"02",x"99",x"ff"),
   603 => (x"f2",x"e7",x"c2",x"87"),
   604 => (x"fd",x"49",x"73",x"1e"),
   605 => (x"86",x"c4",x"87",x"d0"),
   606 => (x"87",x"dc",x"f6",x"26"),
   607 => (x"5c",x"5b",x"5e",x"0e"),
   608 => (x"86",x"f0",x"0e",x"5d"),
   609 => (x"c0",x"59",x"a6",x"d0"),
   610 => (x"cc",x"4b",x"66",x"e4"),
   611 => (x"87",x"ca",x"02",x"66"),
   612 => (x"70",x"80",x"c8",x"48"),
   613 => (x"05",x"bf",x"6e",x"7e"),
   614 => (x"48",x"c0",x"87",x"c5"),
   615 => (x"cc",x"87",x"ec",x"c3"),
   616 => (x"84",x"d0",x"4c",x"66"),
   617 => (x"a6",x"c4",x"49",x"73"),
   618 => (x"c4",x"78",x"6c",x"48"),
   619 => (x"80",x"c4",x"81",x"66"),
   620 => (x"c8",x"78",x"bf",x"6e"),
   621 => (x"c6",x"06",x"a9",x"66"),
   622 => (x"66",x"c4",x"49",x"87"),
   623 => (x"c0",x"4b",x"71",x"89"),
   624 => (x"c4",x"01",x"ab",x"b7"),
   625 => (x"c2",x"c3",x"48",x"87"),
   626 => (x"48",x"66",x"c4",x"87"),
   627 => (x"70",x"98",x"ff",x"c7"),
   628 => (x"c1",x"02",x"6e",x"7e"),
   629 => (x"c0",x"c8",x"87",x"c9"),
   630 => (x"71",x"89",x"6e",x"49"),
   631 => (x"f2",x"e7",x"c2",x"4a"),
   632 => (x"73",x"85",x"6e",x"4d"),
   633 => (x"c1",x"06",x"aa",x"b7"),
   634 => (x"49",x"72",x"4a",x"87"),
   635 => (x"80",x"66",x"c4",x"48"),
   636 => (x"8b",x"72",x"7c",x"70"),
   637 => (x"71",x"8a",x"c1",x"49"),
   638 => (x"87",x"d9",x"02",x"99"),
   639 => (x"48",x"66",x"e0",x"c0"),
   640 => (x"e0",x"c0",x"50",x"15"),
   641 => (x"80",x"c1",x"48",x"66"),
   642 => (x"58",x"a6",x"e4",x"c0"),
   643 => (x"8a",x"c1",x"49",x"72"),
   644 => (x"e7",x"05",x"99",x"71"),
   645 => (x"d0",x"1e",x"c1",x"87"),
   646 => (x"cf",x"f9",x"49",x"66"),
   647 => (x"c0",x"86",x"c4",x"87"),
   648 => (x"c1",x"06",x"ab",x"b7"),
   649 => (x"e0",x"c0",x"87",x"e3"),
   650 => (x"ff",x"c7",x"4d",x"66"),
   651 => (x"c0",x"06",x"ab",x"b7"),
   652 => (x"1e",x"75",x"87",x"e2"),
   653 => (x"fa",x"49",x"66",x"d0"),
   654 => (x"c0",x"c8",x"87",x"cc"),
   655 => (x"c8",x"48",x"6c",x"85"),
   656 => (x"7c",x"70",x"80",x"c0"),
   657 => (x"c1",x"8b",x"c0",x"c8"),
   658 => (x"49",x"66",x"d4",x"1e"),
   659 => (x"c8",x"87",x"dd",x"f8"),
   660 => (x"87",x"ee",x"c0",x"86"),
   661 => (x"1e",x"f2",x"e7",x"c2"),
   662 => (x"f9",x"49",x"66",x"d0"),
   663 => (x"86",x"c4",x"87",x"e8"),
   664 => (x"4a",x"f2",x"e7",x"c2"),
   665 => (x"6c",x"48",x"49",x"73"),
   666 => (x"73",x"7c",x"70",x"80"),
   667 => (x"71",x"8b",x"c1",x"49"),
   668 => (x"87",x"ce",x"02",x"99"),
   669 => (x"c1",x"7d",x"97",x"12"),
   670 => (x"c1",x"49",x"73",x"85"),
   671 => (x"05",x"99",x"71",x"8b"),
   672 => (x"b7",x"c0",x"87",x"f2"),
   673 => (x"e1",x"fe",x"01",x"ab"),
   674 => (x"f0",x"48",x"c1",x"87"),
   675 => (x"87",x"c8",x"f2",x"8e"),
   676 => (x"5c",x"5b",x"5e",x"0e"),
   677 => (x"4b",x"71",x"0e",x"5d"),
   678 => (x"87",x"c7",x"02",x"9b"),
   679 => (x"6d",x"4d",x"a3",x"c8"),
   680 => (x"ff",x"87",x"c5",x"05"),
   681 => (x"87",x"fd",x"c0",x"48"),
   682 => (x"6c",x"4c",x"a3",x"d0"),
   683 => (x"99",x"ff",x"c7",x"49"),
   684 => (x"6c",x"87",x"d8",x"05"),
   685 => (x"c1",x"87",x"c9",x"02"),
   686 => (x"f6",x"49",x"73",x"1e"),
   687 => (x"86",x"c4",x"87",x"ee"),
   688 => (x"1e",x"f2",x"e7",x"c2"),
   689 => (x"fd",x"f7",x"49",x"73"),
   690 => (x"6c",x"86",x"c4",x"87"),
   691 => (x"04",x"aa",x"6d",x"4a"),
   692 => (x"48",x"ff",x"87",x"c4"),
   693 => (x"a2",x"c1",x"87",x"cf"),
   694 => (x"c7",x"49",x"72",x"7c"),
   695 => (x"e7",x"c2",x"99",x"ff"),
   696 => (x"69",x"97",x"81",x"f2"),
   697 => (x"87",x"f0",x"f0",x"48"),
   698 => (x"71",x"1e",x"73",x"1e"),
   699 => (x"c0",x"02",x"9b",x"4b"),
   700 => (x"f4",x"c2",x"87",x"e4"),
   701 => (x"4a",x"73",x"5b",x"df"),
   702 => (x"ef",x"c2",x"8a",x"c2"),
   703 => (x"92",x"49",x"bf",x"f2"),
   704 => (x"bf",x"cb",x"f4",x"c2"),
   705 => (x"c2",x"80",x"72",x"48"),
   706 => (x"71",x"58",x"e3",x"f4"),
   707 => (x"c2",x"30",x"c4",x"48"),
   708 => (x"c0",x"58",x"c2",x"f0"),
   709 => (x"f4",x"c2",x"87",x"ed"),
   710 => (x"f4",x"c2",x"48",x"db"),
   711 => (x"c2",x"78",x"bf",x"cf"),
   712 => (x"c2",x"48",x"df",x"f4"),
   713 => (x"78",x"bf",x"d3",x"f4"),
   714 => (x"bf",x"fa",x"ef",x"c2"),
   715 => (x"c2",x"87",x"c9",x"02"),
   716 => (x"49",x"bf",x"f2",x"ef"),
   717 => (x"87",x"c7",x"31",x"c4"),
   718 => (x"bf",x"d7",x"f4",x"c2"),
   719 => (x"c2",x"31",x"c4",x"49"),
   720 => (x"ef",x"59",x"c2",x"f0"),
   721 => (x"5e",x"0e",x"87",x"d6"),
   722 => (x"71",x"0e",x"5c",x"5b"),
   723 => (x"72",x"4b",x"c0",x"4a"),
   724 => (x"e1",x"c0",x"02",x"9a"),
   725 => (x"49",x"a2",x"da",x"87"),
   726 => (x"c2",x"4b",x"69",x"9f"),
   727 => (x"02",x"bf",x"fa",x"ef"),
   728 => (x"a2",x"d4",x"87",x"cf"),
   729 => (x"49",x"69",x"9f",x"49"),
   730 => (x"ff",x"ff",x"c0",x"4c"),
   731 => (x"c2",x"34",x"d0",x"9c"),
   732 => (x"74",x"4c",x"c0",x"87"),
   733 => (x"49",x"73",x"b3",x"49"),
   734 => (x"ee",x"87",x"ed",x"fd"),
   735 => (x"5e",x"0e",x"87",x"dc"),
   736 => (x"0e",x"5d",x"5c",x"5b"),
   737 => (x"4a",x"71",x"86",x"f4"),
   738 => (x"9a",x"72",x"7e",x"c0"),
   739 => (x"c2",x"87",x"d8",x"02"),
   740 => (x"c0",x"48",x"ee",x"e7"),
   741 => (x"e6",x"e7",x"c2",x"78"),
   742 => (x"df",x"f4",x"c2",x"48"),
   743 => (x"e7",x"c2",x"78",x"bf"),
   744 => (x"f4",x"c2",x"48",x"ea"),
   745 => (x"c2",x"78",x"bf",x"db"),
   746 => (x"c0",x"48",x"cf",x"f0"),
   747 => (x"fe",x"ef",x"c2",x"50"),
   748 => (x"e7",x"c2",x"49",x"bf"),
   749 => (x"71",x"4a",x"bf",x"ee"),
   750 => (x"ca",x"c4",x"03",x"aa"),
   751 => (x"cf",x"49",x"72",x"87"),
   752 => (x"ea",x"c0",x"05",x"99"),
   753 => (x"da",x"f5",x"c0",x"87"),
   754 => (x"e6",x"e7",x"c2",x"48"),
   755 => (x"e7",x"c2",x"78",x"bf"),
   756 => (x"e7",x"c2",x"1e",x"f2"),
   757 => (x"c2",x"49",x"bf",x"e6"),
   758 => (x"c1",x"48",x"e6",x"e7"),
   759 => (x"ff",x"71",x"78",x"a1"),
   760 => (x"c4",x"87",x"f7",x"de"),
   761 => (x"d6",x"f5",x"c0",x"86"),
   762 => (x"f2",x"e7",x"c2",x"48"),
   763 => (x"c0",x"87",x"cc",x"78"),
   764 => (x"48",x"bf",x"d6",x"f5"),
   765 => (x"c0",x"80",x"e0",x"c0"),
   766 => (x"c2",x"58",x"da",x"f5"),
   767 => (x"48",x"bf",x"ee",x"e7"),
   768 => (x"e7",x"c2",x"80",x"c1"),
   769 => (x"56",x"27",x"58",x"f2"),
   770 => (x"bf",x"00",x"00",x"0d"),
   771 => (x"9d",x"4d",x"bf",x"97"),
   772 => (x"87",x"e3",x"c2",x"02"),
   773 => (x"02",x"ad",x"e5",x"c3"),
   774 => (x"c0",x"87",x"dc",x"c2"),
   775 => (x"4b",x"bf",x"d6",x"f5"),
   776 => (x"11",x"49",x"a3",x"cb"),
   777 => (x"05",x"ac",x"cf",x"4c"),
   778 => (x"75",x"87",x"d2",x"c1"),
   779 => (x"c1",x"99",x"df",x"49"),
   780 => (x"c2",x"91",x"cd",x"89"),
   781 => (x"c1",x"81",x"c2",x"f0"),
   782 => (x"51",x"12",x"4a",x"a3"),
   783 => (x"12",x"4a",x"a3",x"c3"),
   784 => (x"4a",x"a3",x"c5",x"51"),
   785 => (x"a3",x"c7",x"51",x"12"),
   786 => (x"c9",x"51",x"12",x"4a"),
   787 => (x"51",x"12",x"4a",x"a3"),
   788 => (x"12",x"4a",x"a3",x"ce"),
   789 => (x"4a",x"a3",x"d0",x"51"),
   790 => (x"a3",x"d2",x"51",x"12"),
   791 => (x"d4",x"51",x"12",x"4a"),
   792 => (x"51",x"12",x"4a",x"a3"),
   793 => (x"12",x"4a",x"a3",x"d6"),
   794 => (x"4a",x"a3",x"d8",x"51"),
   795 => (x"a3",x"dc",x"51",x"12"),
   796 => (x"de",x"51",x"12",x"4a"),
   797 => (x"51",x"12",x"4a",x"a3"),
   798 => (x"fa",x"c0",x"7e",x"c1"),
   799 => (x"c8",x"49",x"74",x"87"),
   800 => (x"eb",x"c0",x"05",x"99"),
   801 => (x"d0",x"49",x"74",x"87"),
   802 => (x"87",x"d1",x"05",x"99"),
   803 => (x"c0",x"02",x"66",x"dc"),
   804 => (x"49",x"73",x"87",x"cb"),
   805 => (x"70",x"0f",x"66",x"dc"),
   806 => (x"d3",x"c0",x"02",x"98"),
   807 => (x"c0",x"05",x"6e",x"87"),
   808 => (x"f0",x"c2",x"87",x"c6"),
   809 => (x"50",x"c0",x"48",x"c2"),
   810 => (x"bf",x"d6",x"f5",x"c0"),
   811 => (x"87",x"e1",x"c2",x"48"),
   812 => (x"48",x"cf",x"f0",x"c2"),
   813 => (x"c2",x"7e",x"50",x"c0"),
   814 => (x"49",x"bf",x"fe",x"ef"),
   815 => (x"bf",x"ee",x"e7",x"c2"),
   816 => (x"04",x"aa",x"71",x"4a"),
   817 => (x"c2",x"87",x"f6",x"fb"),
   818 => (x"05",x"bf",x"df",x"f4"),
   819 => (x"c2",x"87",x"c8",x"c0"),
   820 => (x"02",x"bf",x"fa",x"ef"),
   821 => (x"c2",x"87",x"f8",x"c1"),
   822 => (x"49",x"bf",x"ea",x"e7"),
   823 => (x"70",x"87",x"c1",x"e9"),
   824 => (x"ee",x"e7",x"c2",x"49"),
   825 => (x"48",x"a6",x"c4",x"59"),
   826 => (x"bf",x"ea",x"e7",x"c2"),
   827 => (x"fa",x"ef",x"c2",x"78"),
   828 => (x"d8",x"c0",x"02",x"bf"),
   829 => (x"49",x"66",x"c4",x"87"),
   830 => (x"ff",x"ff",x"ff",x"cf"),
   831 => (x"02",x"a9",x"99",x"f8"),
   832 => (x"c0",x"87",x"c5",x"c0"),
   833 => (x"87",x"e1",x"c0",x"4c"),
   834 => (x"dc",x"c0",x"4c",x"c1"),
   835 => (x"49",x"66",x"c4",x"87"),
   836 => (x"99",x"f8",x"ff",x"cf"),
   837 => (x"c8",x"c0",x"02",x"a9"),
   838 => (x"48",x"a6",x"c8",x"87"),
   839 => (x"c5",x"c0",x"78",x"c0"),
   840 => (x"48",x"a6",x"c8",x"87"),
   841 => (x"66",x"c8",x"78",x"c1"),
   842 => (x"05",x"9c",x"74",x"4c"),
   843 => (x"c4",x"87",x"e0",x"c0"),
   844 => (x"89",x"c2",x"49",x"66"),
   845 => (x"bf",x"f2",x"ef",x"c2"),
   846 => (x"f4",x"c2",x"91",x"4a"),
   847 => (x"c2",x"4a",x"bf",x"cb"),
   848 => (x"72",x"48",x"e6",x"e7"),
   849 => (x"e7",x"c2",x"78",x"a1"),
   850 => (x"78",x"c0",x"48",x"ee"),
   851 => (x"c0",x"87",x"de",x"f9"),
   852 => (x"e7",x"8e",x"f4",x"48"),
   853 => (x"00",x"00",x"87",x"c2"),
   854 => (x"ff",x"ff",x"00",x"00"),
   855 => (x"0d",x"66",x"ff",x"ff"),
   856 => (x"0d",x"6f",x"00",x"00"),
   857 => (x"41",x"46",x"00",x"00"),
   858 => (x"20",x"32",x"33",x"54"),
   859 => (x"46",x"00",x"20",x"20"),
   860 => (x"36",x"31",x"54",x"41"),
   861 => (x"00",x"20",x"20",x"20"),
   862 => (x"e4",x"f4",x"c2",x"1e"),
   863 => (x"a8",x"dd",x"48",x"bf"),
   864 => (x"c1",x"87",x"c9",x"05"),
   865 => (x"70",x"87",x"e3",x"c2"),
   866 => (x"87",x"c8",x"4a",x"49"),
   867 => (x"c3",x"48",x"d4",x"ff"),
   868 => (x"4a",x"68",x"78",x"ff"),
   869 => (x"4f",x"26",x"48",x"72"),
   870 => (x"e4",x"f4",x"c2",x"1e"),
   871 => (x"a8",x"dd",x"48",x"bf"),
   872 => (x"c1",x"87",x"c6",x"05"),
   873 => (x"d9",x"87",x"ef",x"c1"),
   874 => (x"48",x"d4",x"ff",x"87"),
   875 => (x"ff",x"78",x"ff",x"c3"),
   876 => (x"e1",x"c0",x"48",x"d0"),
   877 => (x"48",x"d4",x"ff",x"78"),
   878 => (x"f4",x"c2",x"78",x"d4"),
   879 => (x"d4",x"ff",x"48",x"e3"),
   880 => (x"4f",x"26",x"50",x"bf"),
   881 => (x"48",x"d0",x"ff",x"1e"),
   882 => (x"26",x"78",x"e0",x"c0"),
   883 => (x"e7",x"fe",x"1e",x"4f"),
   884 => (x"99",x"49",x"70",x"87"),
   885 => (x"c0",x"87",x"c6",x"02"),
   886 => (x"f1",x"05",x"a9",x"fb"),
   887 => (x"26",x"48",x"71",x"87"),
   888 => (x"5b",x"5e",x"0e",x"4f"),
   889 => (x"4b",x"71",x"0e",x"5c"),
   890 => (x"cb",x"fe",x"4c",x"c0"),
   891 => (x"99",x"49",x"70",x"87"),
   892 => (x"87",x"f9",x"c0",x"02"),
   893 => (x"02",x"a9",x"ec",x"c0"),
   894 => (x"c0",x"87",x"f2",x"c0"),
   895 => (x"c0",x"02",x"a9",x"fb"),
   896 => (x"66",x"cc",x"87",x"eb"),
   897 => (x"c7",x"03",x"ac",x"b7"),
   898 => (x"02",x"66",x"d0",x"87"),
   899 => (x"53",x"71",x"87",x"c2"),
   900 => (x"c2",x"02",x"99",x"71"),
   901 => (x"fd",x"84",x"c1",x"87"),
   902 => (x"49",x"70",x"87",x"de"),
   903 => (x"87",x"cd",x"02",x"99"),
   904 => (x"02",x"a9",x"ec",x"c0"),
   905 => (x"fb",x"c0",x"87",x"c7"),
   906 => (x"d5",x"ff",x"05",x"a9"),
   907 => (x"02",x"66",x"d0",x"87"),
   908 => (x"97",x"c0",x"87",x"c3"),
   909 => (x"a9",x"ec",x"c0",x"7b"),
   910 => (x"74",x"87",x"c4",x"05"),
   911 => (x"74",x"87",x"c5",x"4a"),
   912 => (x"8a",x"0a",x"c0",x"4a"),
   913 => (x"87",x"c2",x"48",x"72"),
   914 => (x"4c",x"26",x"4d",x"26"),
   915 => (x"4f",x"26",x"4b",x"26"),
   916 => (x"87",x"e4",x"fc",x"1e"),
   917 => (x"f0",x"c0",x"49",x"70"),
   918 => (x"ca",x"04",x"a9",x"b7"),
   919 => (x"b7",x"f9",x"c0",x"87"),
   920 => (x"87",x"c3",x"01",x"a9"),
   921 => (x"c1",x"89",x"f0",x"c0"),
   922 => (x"04",x"a9",x"b7",x"c1"),
   923 => (x"da",x"c1",x"87",x"ca"),
   924 => (x"c3",x"01",x"a9",x"b7"),
   925 => (x"89",x"f7",x"c0",x"87"),
   926 => (x"4f",x"26",x"48",x"71"),
   927 => (x"5c",x"5b",x"5e",x"0e"),
   928 => (x"fc",x"4c",x"71",x"0e"),
   929 => (x"1e",x"c1",x"87",x"d2"),
   930 => (x"74",x"1e",x"66",x"d0"),
   931 => (x"87",x"d1",x"fd",x"49"),
   932 => (x"4b",x"70",x"86",x"c8"),
   933 => (x"c0",x"87",x"ed",x"fc"),
   934 => (x"c2",x"03",x"ab",x"b7"),
   935 => (x"cc",x"8b",x"0b",x"87"),
   936 => (x"03",x"ab",x"b7",x"66"),
   937 => (x"a3",x"74",x"87",x"cf"),
   938 => (x"c0",x"83",x"c1",x"49"),
   939 => (x"66",x"cc",x"51",x"e0"),
   940 => (x"f1",x"04",x"ab",x"b7"),
   941 => (x"49",x"a3",x"74",x"87"),
   942 => (x"cd",x"fe",x"51",x"c0"),
   943 => (x"5b",x"5e",x"0e",x"87"),
   944 => (x"4a",x"71",x"0e",x"5c"),
   945 => (x"72",x"4c",x"d4",x"ff"),
   946 => (x"87",x"e9",x"c0",x"49"),
   947 => (x"02",x"9b",x"4b",x"70"),
   948 => (x"8b",x"c1",x"87",x"c2"),
   949 => (x"c5",x"48",x"d0",x"ff"),
   950 => (x"7c",x"d5",x"c1",x"78"),
   951 => (x"31",x"c6",x"49",x"73"),
   952 => (x"97",x"d7",x"e7",x"c1"),
   953 => (x"71",x"48",x"4a",x"bf"),
   954 => (x"ff",x"7c",x"70",x"b0"),
   955 => (x"78",x"c4",x"48",x"d0"),
   956 => (x"d5",x"fd",x"48",x"73"),
   957 => (x"5b",x"5e",x"0e",x"87"),
   958 => (x"f4",x"0e",x"5d",x"5c"),
   959 => (x"c4",x"4c",x"71",x"86"),
   960 => (x"78",x"c0",x"48",x"a6"),
   961 => (x"6e",x"7e",x"a4",x"c8"),
   962 => (x"c1",x"49",x"bf",x"97"),
   963 => (x"dd",x"05",x"a9",x"c1"),
   964 => (x"49",x"a4",x"c9",x"87"),
   965 => (x"c1",x"49",x"69",x"97"),
   966 => (x"d1",x"05",x"a9",x"d2"),
   967 => (x"49",x"a4",x"ca",x"87"),
   968 => (x"c1",x"49",x"69",x"97"),
   969 => (x"c5",x"05",x"a9",x"c3"),
   970 => (x"c2",x"48",x"df",x"87"),
   971 => (x"e7",x"f9",x"87",x"e1"),
   972 => (x"c0",x"4b",x"c0",x"87"),
   973 => (x"bf",x"97",x"d4",x"ff"),
   974 => (x"04",x"a9",x"c0",x"49"),
   975 => (x"cc",x"fa",x"87",x"cf"),
   976 => (x"c0",x"83",x"c1",x"87"),
   977 => (x"bf",x"97",x"d4",x"ff"),
   978 => (x"f1",x"06",x"ab",x"49"),
   979 => (x"d4",x"ff",x"c0",x"87"),
   980 => (x"cf",x"02",x"bf",x"97"),
   981 => (x"87",x"e0",x"f8",x"87"),
   982 => (x"02",x"99",x"49",x"70"),
   983 => (x"ec",x"c0",x"87",x"c6"),
   984 => (x"87",x"f1",x"05",x"a9"),
   985 => (x"cf",x"f8",x"4b",x"c0"),
   986 => (x"f8",x"4d",x"70",x"87"),
   987 => (x"a6",x"cc",x"87",x"ca"),
   988 => (x"87",x"c4",x"f8",x"58"),
   989 => (x"83",x"c1",x"4a",x"70"),
   990 => (x"49",x"bf",x"97",x"6e"),
   991 => (x"87",x"c7",x"02",x"ad"),
   992 => (x"05",x"ad",x"ff",x"c0"),
   993 => (x"c9",x"87",x"ea",x"c0"),
   994 => (x"69",x"97",x"49",x"a4"),
   995 => (x"a9",x"66",x"c8",x"49"),
   996 => (x"48",x"87",x"c7",x"02"),
   997 => (x"05",x"a8",x"ff",x"c0"),
   998 => (x"a4",x"ca",x"87",x"d7"),
   999 => (x"49",x"69",x"97",x"49"),
  1000 => (x"87",x"c6",x"02",x"aa"),
  1001 => (x"05",x"aa",x"ff",x"c0"),
  1002 => (x"a6",x"c4",x"87",x"c7"),
  1003 => (x"d3",x"78",x"c1",x"48"),
  1004 => (x"ad",x"ec",x"c0",x"87"),
  1005 => (x"c0",x"87",x"c6",x"02"),
  1006 => (x"c7",x"05",x"ad",x"fb"),
  1007 => (x"c4",x"4b",x"c0",x"87"),
  1008 => (x"78",x"c1",x"48",x"a6"),
  1009 => (x"fe",x"02",x"66",x"c4"),
  1010 => (x"f7",x"f7",x"87",x"dc"),
  1011 => (x"f4",x"48",x"73",x"87"),
  1012 => (x"87",x"f4",x"f9",x"8e"),
  1013 => (x"5b",x"5e",x"0e",x"00"),
  1014 => (x"1e",x"0e",x"5d",x"5c"),
  1015 => (x"d4",x"ff",x"4d",x"71"),
  1016 => (x"c2",x"1e",x"75",x"4b"),
  1017 => (x"e0",x"49",x"e8",x"f4"),
  1018 => (x"86",x"c4",x"87",x"c7"),
  1019 => (x"c4",x"02",x"98",x"70"),
  1020 => (x"f4",x"c2",x"87",x"c8"),
  1021 => (x"75",x"4c",x"bf",x"f0"),
  1022 => (x"87",x"c1",x"fb",x"49"),
  1023 => (x"c0",x"05",x"a8",x"de"),
  1024 => (x"49",x"75",x"87",x"eb"),
  1025 => (x"87",x"c0",x"f6",x"c0"),
  1026 => (x"db",x"02",x"98",x"70"),
  1027 => (x"cc",x"f9",x"c2",x"87"),
  1028 => (x"e1",x"c0",x"1e",x"bf"),
  1029 => (x"cf",x"f3",x"c0",x"49"),
  1030 => (x"c1",x"86",x"c4",x"87"),
  1031 => (x"c0",x"48",x"d7",x"e7"),
  1032 => (x"d8",x"f9",x"c2",x"50"),
  1033 => (x"87",x"ed",x"fe",x"49"),
  1034 => (x"cf",x"c3",x"48",x"c1"),
  1035 => (x"48",x"d0",x"ff",x"87"),
  1036 => (x"d6",x"c1",x"78",x"c5"),
  1037 => (x"75",x"4a",x"c0",x"7b"),
  1038 => (x"7b",x"11",x"49",x"a2"),
  1039 => (x"b7",x"cb",x"82",x"c1"),
  1040 => (x"87",x"f3",x"04",x"aa"),
  1041 => (x"ff",x"c3",x"4a",x"cc"),
  1042 => (x"c0",x"82",x"c1",x"7b"),
  1043 => (x"04",x"aa",x"b7",x"e0"),
  1044 => (x"d0",x"ff",x"87",x"f4"),
  1045 => (x"c3",x"78",x"c4",x"48"),
  1046 => (x"78",x"c5",x"7b",x"ff"),
  1047 => (x"c1",x"7b",x"d3",x"c1"),
  1048 => (x"74",x"78",x"c4",x"7b"),
  1049 => (x"c0",x"c2",x"02",x"9c"),
  1050 => (x"f2",x"e7",x"c2",x"87"),
  1051 => (x"4d",x"c0",x"c8",x"7e"),
  1052 => (x"ac",x"b7",x"c0",x"8c"),
  1053 => (x"c8",x"87",x"c6",x"03"),
  1054 => (x"c0",x"4d",x"a4",x"c0"),
  1055 => (x"ad",x"c0",x"c8",x"4c"),
  1056 => (x"c2",x"87",x"dc",x"05"),
  1057 => (x"bf",x"97",x"e3",x"f4"),
  1058 => (x"02",x"99",x"d0",x"49"),
  1059 => (x"1e",x"c0",x"87",x"d1"),
  1060 => (x"49",x"e8",x"f4",x"c2"),
  1061 => (x"c4",x"87",x"ef",x"e0"),
  1062 => (x"4a",x"49",x"70",x"86"),
  1063 => (x"c2",x"87",x"ee",x"c0"),
  1064 => (x"c2",x"1e",x"f2",x"e7"),
  1065 => (x"e0",x"49",x"e8",x"f4"),
  1066 => (x"86",x"c4",x"87",x"dc"),
  1067 => (x"ff",x"4a",x"49",x"70"),
  1068 => (x"c5",x"c8",x"48",x"d0"),
  1069 => (x"7b",x"d4",x"c1",x"78"),
  1070 => (x"7b",x"bf",x"97",x"6e"),
  1071 => (x"80",x"c1",x"48",x"6e"),
  1072 => (x"8d",x"c1",x"7e",x"70"),
  1073 => (x"87",x"f0",x"ff",x"05"),
  1074 => (x"c4",x"48",x"d0",x"ff"),
  1075 => (x"05",x"9a",x"72",x"78"),
  1076 => (x"48",x"c0",x"87",x"c5"),
  1077 => (x"c1",x"87",x"e5",x"c0"),
  1078 => (x"e8",x"f4",x"c2",x"1e"),
  1079 => (x"cb",x"de",x"ff",x"49"),
  1080 => (x"74",x"86",x"c4",x"87"),
  1081 => (x"c0",x"fe",x"05",x"9c"),
  1082 => (x"48",x"d0",x"ff",x"87"),
  1083 => (x"d3",x"c1",x"78",x"c5"),
  1084 => (x"c4",x"7b",x"c0",x"7b"),
  1085 => (x"c0",x"48",x"c1",x"78"),
  1086 => (x"48",x"c0",x"87",x"c2"),
  1087 => (x"26",x"4d",x"26",x"26"),
  1088 => (x"26",x"4b",x"26",x"4c"),
  1089 => (x"5b",x"5e",x"0e",x"4f"),
  1090 => (x"1e",x"0e",x"5d",x"5c"),
  1091 => (x"4c",x"c0",x"4b",x"71"),
  1092 => (x"c0",x"04",x"ab",x"4d"),
  1093 => (x"fb",x"c0",x"87",x"e8"),
  1094 => (x"9d",x"75",x"1e",x"f5"),
  1095 => (x"c0",x"87",x"c4",x"02"),
  1096 => (x"c1",x"87",x"c2",x"4a"),
  1097 => (x"e9",x"49",x"72",x"4a"),
  1098 => (x"86",x"c4",x"87",x"d4"),
  1099 => (x"84",x"c1",x"7e",x"70"),
  1100 => (x"87",x"c2",x"05",x"6e"),
  1101 => (x"85",x"c1",x"4c",x"73"),
  1102 => (x"ff",x"06",x"ac",x"73"),
  1103 => (x"48",x"6e",x"87",x"d8"),
  1104 => (x"87",x"f9",x"fe",x"26"),
  1105 => (x"c4",x"4a",x"71",x"1e"),
  1106 => (x"87",x"c5",x"05",x"66"),
  1107 => (x"c4",x"fa",x"49",x"72"),
  1108 => (x"0e",x"4f",x"26",x"87"),
  1109 => (x"5d",x"5c",x"5b",x"5e"),
  1110 => (x"4c",x"71",x"1e",x"0e"),
  1111 => (x"c2",x"91",x"de",x"49"),
  1112 => (x"71",x"4d",x"d0",x"f5"),
  1113 => (x"02",x"6d",x"97",x"85"),
  1114 => (x"c2",x"87",x"dc",x"c1"),
  1115 => (x"4a",x"bf",x"fc",x"f4"),
  1116 => (x"49",x"72",x"82",x"74"),
  1117 => (x"70",x"87",x"ce",x"fe"),
  1118 => (x"c0",x"02",x"6e",x"7e"),
  1119 => (x"f5",x"c2",x"87",x"f2"),
  1120 => (x"4a",x"6e",x"4b",x"c4"),
  1121 => (x"fc",x"fe",x"49",x"cb"),
  1122 => (x"4b",x"74",x"87",x"de"),
  1123 => (x"e7",x"c1",x"93",x"cb"),
  1124 => (x"83",x"c4",x"83",x"e7"),
  1125 => (x"7b",x"cb",x"c7",x"c1"),
  1126 => (x"cb",x"c1",x"49",x"74"),
  1127 => (x"7b",x"75",x"87",x"d7"),
  1128 => (x"97",x"d8",x"e7",x"c1"),
  1129 => (x"c2",x"1e",x"49",x"bf"),
  1130 => (x"fe",x"49",x"c4",x"f5"),
  1131 => (x"86",x"c4",x"87",x"d6"),
  1132 => (x"ca",x"c1",x"49",x"74"),
  1133 => (x"49",x"c0",x"87",x"ff"),
  1134 => (x"87",x"de",x"cc",x"c1"),
  1135 => (x"48",x"e4",x"f4",x"c2"),
  1136 => (x"49",x"c1",x"78",x"c0"),
  1137 => (x"26",x"87",x"cf",x"dd"),
  1138 => (x"4c",x"87",x"f2",x"fc"),
  1139 => (x"69",x"64",x"61",x"6f"),
  1140 => (x"2e",x"2e",x"67",x"6e"),
  1141 => (x"5e",x"0e",x"00",x"2e"),
  1142 => (x"71",x"0e",x"5c",x"5b"),
  1143 => (x"f4",x"c2",x"4a",x"4b"),
  1144 => (x"72",x"82",x"bf",x"fc"),
  1145 => (x"87",x"dd",x"fc",x"49"),
  1146 => (x"02",x"9c",x"4c",x"70"),
  1147 => (x"e5",x"49",x"87",x"c4"),
  1148 => (x"f4",x"c2",x"87",x"d4"),
  1149 => (x"78",x"c0",x"48",x"fc"),
  1150 => (x"d9",x"dc",x"49",x"c1"),
  1151 => (x"87",x"ff",x"fb",x"87"),
  1152 => (x"5c",x"5b",x"5e",x"0e"),
  1153 => (x"86",x"f4",x"0e",x"5d"),
  1154 => (x"4d",x"f2",x"e7",x"c2"),
  1155 => (x"a6",x"c4",x"4c",x"c0"),
  1156 => (x"c2",x"78",x"c0",x"48"),
  1157 => (x"49",x"bf",x"fc",x"f4"),
  1158 => (x"c1",x"06",x"a9",x"c0"),
  1159 => (x"e7",x"c2",x"87",x"c1"),
  1160 => (x"02",x"98",x"48",x"f2"),
  1161 => (x"c0",x"87",x"f8",x"c0"),
  1162 => (x"c8",x"1e",x"f5",x"fb"),
  1163 => (x"87",x"c7",x"02",x"66"),
  1164 => (x"c0",x"48",x"a6",x"c4"),
  1165 => (x"c4",x"87",x"c5",x"78"),
  1166 => (x"78",x"c1",x"48",x"a6"),
  1167 => (x"e4",x"49",x"66",x"c4"),
  1168 => (x"86",x"c4",x"87",x"fc"),
  1169 => (x"84",x"c1",x"4d",x"70"),
  1170 => (x"c1",x"48",x"66",x"c4"),
  1171 => (x"58",x"a6",x"c8",x"80"),
  1172 => (x"bf",x"fc",x"f4",x"c2"),
  1173 => (x"c6",x"03",x"ac",x"49"),
  1174 => (x"05",x"9d",x"75",x"87"),
  1175 => (x"c0",x"87",x"c8",x"ff"),
  1176 => (x"02",x"9d",x"75",x"4c"),
  1177 => (x"c0",x"87",x"e0",x"c3"),
  1178 => (x"c8",x"1e",x"f5",x"fb"),
  1179 => (x"87",x"c7",x"02",x"66"),
  1180 => (x"c0",x"48",x"a6",x"cc"),
  1181 => (x"cc",x"87",x"c5",x"78"),
  1182 => (x"78",x"c1",x"48",x"a6"),
  1183 => (x"e3",x"49",x"66",x"cc"),
  1184 => (x"86",x"c4",x"87",x"fc"),
  1185 => (x"02",x"6e",x"7e",x"70"),
  1186 => (x"6e",x"87",x"e9",x"c2"),
  1187 => (x"97",x"81",x"cb",x"49"),
  1188 => (x"99",x"d0",x"49",x"69"),
  1189 => (x"87",x"d6",x"c1",x"02"),
  1190 => (x"4a",x"d6",x"c7",x"c1"),
  1191 => (x"91",x"cb",x"49",x"74"),
  1192 => (x"81",x"e7",x"e7",x"c1"),
  1193 => (x"81",x"c8",x"79",x"72"),
  1194 => (x"74",x"51",x"ff",x"c3"),
  1195 => (x"c2",x"91",x"de",x"49"),
  1196 => (x"71",x"4d",x"d0",x"f5"),
  1197 => (x"97",x"c1",x"c2",x"85"),
  1198 => (x"49",x"a5",x"c1",x"7d"),
  1199 => (x"c2",x"51",x"e0",x"c0"),
  1200 => (x"bf",x"97",x"c2",x"f0"),
  1201 => (x"c1",x"87",x"d2",x"02"),
  1202 => (x"4b",x"a5",x"c2",x"84"),
  1203 => (x"4a",x"c2",x"f0",x"c2"),
  1204 => (x"f7",x"fe",x"49",x"db"),
  1205 => (x"db",x"c1",x"87",x"d2"),
  1206 => (x"49",x"a5",x"cd",x"87"),
  1207 => (x"84",x"c1",x"51",x"c0"),
  1208 => (x"6e",x"4b",x"a5",x"c2"),
  1209 => (x"fe",x"49",x"cb",x"4a"),
  1210 => (x"c1",x"87",x"fd",x"f6"),
  1211 => (x"c5",x"c1",x"87",x"c6"),
  1212 => (x"49",x"74",x"4a",x"d3"),
  1213 => (x"e7",x"c1",x"91",x"cb"),
  1214 => (x"79",x"72",x"81",x"e7"),
  1215 => (x"97",x"c2",x"f0",x"c2"),
  1216 => (x"87",x"d8",x"02",x"bf"),
  1217 => (x"91",x"de",x"49",x"74"),
  1218 => (x"f5",x"c2",x"84",x"c1"),
  1219 => (x"83",x"71",x"4b",x"d0"),
  1220 => (x"4a",x"c2",x"f0",x"c2"),
  1221 => (x"f6",x"fe",x"49",x"dd"),
  1222 => (x"87",x"d8",x"87",x"ce"),
  1223 => (x"93",x"de",x"4b",x"74"),
  1224 => (x"83",x"d0",x"f5",x"c2"),
  1225 => (x"c0",x"49",x"a3",x"cb"),
  1226 => (x"73",x"84",x"c1",x"51"),
  1227 => (x"49",x"cb",x"4a",x"6e"),
  1228 => (x"87",x"f4",x"f5",x"fe"),
  1229 => (x"c1",x"48",x"66",x"c4"),
  1230 => (x"58",x"a6",x"c8",x"80"),
  1231 => (x"c0",x"03",x"ac",x"c7"),
  1232 => (x"05",x"6e",x"87",x"c5"),
  1233 => (x"74",x"87",x"e0",x"fc"),
  1234 => (x"f6",x"8e",x"f4",x"48"),
  1235 => (x"73",x"1e",x"87",x"ef"),
  1236 => (x"49",x"4b",x"71",x"1e"),
  1237 => (x"e7",x"c1",x"91",x"cb"),
  1238 => (x"a1",x"c8",x"81",x"e7"),
  1239 => (x"d7",x"e7",x"c1",x"4a"),
  1240 => (x"c9",x"50",x"12",x"48"),
  1241 => (x"ff",x"c0",x"4a",x"a1"),
  1242 => (x"50",x"12",x"48",x"d4"),
  1243 => (x"e7",x"c1",x"81",x"ca"),
  1244 => (x"50",x"11",x"48",x"d8"),
  1245 => (x"97",x"d8",x"e7",x"c1"),
  1246 => (x"c0",x"1e",x"49",x"bf"),
  1247 => (x"87",x"c4",x"f7",x"49"),
  1248 => (x"48",x"e4",x"f4",x"c2"),
  1249 => (x"49",x"c1",x"78",x"de"),
  1250 => (x"26",x"87",x"cb",x"d6"),
  1251 => (x"1e",x"87",x"f2",x"f5"),
  1252 => (x"cb",x"49",x"4a",x"71"),
  1253 => (x"e7",x"e7",x"c1",x"91"),
  1254 => (x"11",x"81",x"c8",x"81"),
  1255 => (x"e8",x"f4",x"c2",x"48"),
  1256 => (x"fc",x"f4",x"c2",x"58"),
  1257 => (x"c1",x"78",x"c0",x"48"),
  1258 => (x"87",x"ea",x"d5",x"49"),
  1259 => (x"c0",x"1e",x"4f",x"26"),
  1260 => (x"e5",x"c4",x"c1",x"49"),
  1261 => (x"1e",x"4f",x"26",x"87"),
  1262 => (x"d2",x"02",x"99",x"71"),
  1263 => (x"fc",x"e8",x"c1",x"87"),
  1264 => (x"f7",x"50",x"c0",x"48"),
  1265 => (x"cf",x"ce",x"c1",x"80"),
  1266 => (x"e0",x"e7",x"c1",x"40"),
  1267 => (x"c1",x"87",x"ce",x"78"),
  1268 => (x"c1",x"48",x"f8",x"e8"),
  1269 => (x"fc",x"78",x"d9",x"e7"),
  1270 => (x"ee",x"ce",x"c1",x"80"),
  1271 => (x"0e",x"4f",x"26",x"78"),
  1272 => (x"0e",x"5c",x"5b",x"5e"),
  1273 => (x"cb",x"4a",x"4c",x"71"),
  1274 => (x"e7",x"e7",x"c1",x"92"),
  1275 => (x"49",x"a2",x"c8",x"82"),
  1276 => (x"97",x"4b",x"a2",x"c9"),
  1277 => (x"97",x"1e",x"4b",x"6b"),
  1278 => (x"ca",x"1e",x"49",x"69"),
  1279 => (x"c0",x"49",x"12",x"82"),
  1280 => (x"c0",x"87",x"c5",x"e5"),
  1281 => (x"87",x"ce",x"d4",x"49"),
  1282 => (x"c1",x"c1",x"49",x"74"),
  1283 => (x"8e",x"f8",x"87",x"e7"),
  1284 => (x"1e",x"87",x"ec",x"f3"),
  1285 => (x"4b",x"71",x"1e",x"73"),
  1286 => (x"87",x"c3",x"ff",x"49"),
  1287 => (x"fe",x"fe",x"49",x"73"),
  1288 => (x"87",x"dd",x"f3",x"87"),
  1289 => (x"71",x"1e",x"73",x"1e"),
  1290 => (x"4a",x"a3",x"c6",x"4b"),
  1291 => (x"c1",x"87",x"db",x"02"),
  1292 => (x"87",x"d6",x"02",x"8a"),
  1293 => (x"da",x"c1",x"02",x"8a"),
  1294 => (x"c0",x"02",x"8a",x"87"),
  1295 => (x"02",x"8a",x"87",x"fc"),
  1296 => (x"8a",x"87",x"e1",x"c0"),
  1297 => (x"c1",x"87",x"cb",x"02"),
  1298 => (x"49",x"c7",x"87",x"db"),
  1299 => (x"c1",x"87",x"c0",x"fd"),
  1300 => (x"f4",x"c2",x"87",x"de"),
  1301 => (x"c1",x"02",x"bf",x"fc"),
  1302 => (x"c1",x"48",x"87",x"cb"),
  1303 => (x"c0",x"f5",x"c2",x"88"),
  1304 => (x"87",x"c1",x"c1",x"58"),
  1305 => (x"bf",x"c0",x"f5",x"c2"),
  1306 => (x"87",x"f9",x"c0",x"02"),
  1307 => (x"bf",x"fc",x"f4",x"c2"),
  1308 => (x"c2",x"80",x"c1",x"48"),
  1309 => (x"c0",x"58",x"c0",x"f5"),
  1310 => (x"f4",x"c2",x"87",x"eb"),
  1311 => (x"c6",x"49",x"bf",x"fc"),
  1312 => (x"c0",x"f5",x"c2",x"89"),
  1313 => (x"a9",x"b7",x"c0",x"59"),
  1314 => (x"c2",x"87",x"da",x"03"),
  1315 => (x"c0",x"48",x"fc",x"f4"),
  1316 => (x"c2",x"87",x"d2",x"78"),
  1317 => (x"02",x"bf",x"c0",x"f5"),
  1318 => (x"f4",x"c2",x"87",x"cb"),
  1319 => (x"c6",x"48",x"bf",x"fc"),
  1320 => (x"c0",x"f5",x"c2",x"80"),
  1321 => (x"d1",x"49",x"c0",x"58"),
  1322 => (x"49",x"73",x"87",x"ec"),
  1323 => (x"87",x"c5",x"ff",x"c0"),
  1324 => (x"1e",x"87",x"ce",x"f1"),
  1325 => (x"4b",x"71",x"1e",x"73"),
  1326 => (x"48",x"e4",x"f4",x"c2"),
  1327 => (x"49",x"c0",x"78",x"dd"),
  1328 => (x"73",x"87",x"d3",x"d1"),
  1329 => (x"ec",x"fe",x"c0",x"49"),
  1330 => (x"87",x"f5",x"f0",x"87"),
  1331 => (x"5c",x"5b",x"5e",x"0e"),
  1332 => (x"cc",x"4c",x"71",x"0e"),
  1333 => (x"4b",x"74",x"1e",x"66"),
  1334 => (x"e7",x"c1",x"93",x"cb"),
  1335 => (x"a3",x"c4",x"83",x"e7"),
  1336 => (x"fe",x"49",x"6a",x"4a"),
  1337 => (x"c1",x"87",x"d1",x"ef"),
  1338 => (x"c8",x"7b",x"ce",x"cd"),
  1339 => (x"66",x"d4",x"49",x"a3"),
  1340 => (x"49",x"a3",x"c9",x"51"),
  1341 => (x"ca",x"51",x"66",x"d8"),
  1342 => (x"66",x"dc",x"49",x"a3"),
  1343 => (x"fe",x"ef",x"26",x"51"),
  1344 => (x"5b",x"5e",x"0e",x"87"),
  1345 => (x"ff",x"0e",x"5d",x"5c"),
  1346 => (x"a6",x"dc",x"86",x"cc"),
  1347 => (x"48",x"a6",x"c8",x"59"),
  1348 => (x"80",x"c4",x"78",x"c0"),
  1349 => (x"78",x"66",x"c8",x"c1"),
  1350 => (x"78",x"c1",x"80",x"c4"),
  1351 => (x"78",x"c1",x"80",x"c4"),
  1352 => (x"48",x"c0",x"f5",x"c2"),
  1353 => (x"f4",x"c2",x"78",x"c1"),
  1354 => (x"de",x"48",x"bf",x"e4"),
  1355 => (x"87",x"cb",x"05",x"a8"),
  1356 => (x"70",x"87",x"cd",x"f3"),
  1357 => (x"59",x"a6",x"cc",x"49"),
  1358 => (x"e1",x"87",x"d6",x"ce"),
  1359 => (x"cc",x"e2",x"87",x"da"),
  1360 => (x"87",x"f4",x"e0",x"87"),
  1361 => (x"fb",x"c0",x"4c",x"70"),
  1362 => (x"d8",x"c1",x"02",x"ac"),
  1363 => (x"05",x"66",x"d8",x"87"),
  1364 => (x"c0",x"87",x"ca",x"c1"),
  1365 => (x"1e",x"c1",x"1e",x"1e"),
  1366 => (x"1e",x"ca",x"e9",x"c1"),
  1367 => (x"eb",x"fd",x"49",x"c0"),
  1368 => (x"c0",x"86",x"d0",x"87"),
  1369 => (x"d9",x"02",x"ac",x"fb"),
  1370 => (x"66",x"c4",x"c1",x"87"),
  1371 => (x"6a",x"82",x"c4",x"4a"),
  1372 => (x"74",x"81",x"c7",x"49"),
  1373 => (x"d8",x"1e",x"c1",x"51"),
  1374 => (x"c8",x"49",x"6a",x"1e"),
  1375 => (x"87",x"e1",x"e1",x"81"),
  1376 => (x"c8",x"c1",x"86",x"c8"),
  1377 => (x"a8",x"c0",x"48",x"66"),
  1378 => (x"c8",x"87",x"c7",x"01"),
  1379 => (x"78",x"c1",x"48",x"a6"),
  1380 => (x"c8",x"c1",x"87",x"ce"),
  1381 => (x"88",x"c1",x"48",x"66"),
  1382 => (x"c3",x"58",x"a6",x"d0"),
  1383 => (x"87",x"ed",x"e0",x"87"),
  1384 => (x"c2",x"48",x"a6",x"d0"),
  1385 => (x"02",x"9c",x"74",x"78"),
  1386 => (x"c8",x"87",x"e2",x"cc"),
  1387 => (x"cc",x"c1",x"48",x"66"),
  1388 => (x"cc",x"03",x"a8",x"66"),
  1389 => (x"a6",x"c4",x"87",x"d7"),
  1390 => (x"d8",x"78",x"c0",x"48"),
  1391 => (x"ff",x"78",x"c0",x"80"),
  1392 => (x"70",x"87",x"f5",x"de"),
  1393 => (x"48",x"66",x"d8",x"4c"),
  1394 => (x"c6",x"05",x"a8",x"dd"),
  1395 => (x"48",x"a6",x"dc",x"87"),
  1396 => (x"c1",x"78",x"66",x"d8"),
  1397 => (x"c0",x"05",x"ac",x"d0"),
  1398 => (x"de",x"ff",x"87",x"eb"),
  1399 => (x"de",x"ff",x"87",x"da"),
  1400 => (x"4c",x"70",x"87",x"d6"),
  1401 => (x"05",x"ac",x"ec",x"c0"),
  1402 => (x"df",x"ff",x"87",x"c6"),
  1403 => (x"4c",x"70",x"87",x"df"),
  1404 => (x"05",x"ac",x"d0",x"c1"),
  1405 => (x"66",x"d4",x"87",x"c8"),
  1406 => (x"d8",x"80",x"c1",x"48"),
  1407 => (x"d0",x"c1",x"58",x"a6"),
  1408 => (x"d5",x"ff",x"02",x"ac"),
  1409 => (x"a6",x"e0",x"c0",x"87"),
  1410 => (x"78",x"66",x"d8",x"48"),
  1411 => (x"c0",x"48",x"66",x"dc"),
  1412 => (x"05",x"a8",x"66",x"e0"),
  1413 => (x"c0",x"87",x"c8",x"ca"),
  1414 => (x"c0",x"48",x"a6",x"e4"),
  1415 => (x"c0",x"80",x"c4",x"78"),
  1416 => (x"c0",x"4d",x"74",x"78"),
  1417 => (x"c9",x"02",x"8d",x"fb"),
  1418 => (x"8d",x"c9",x"87",x"ce"),
  1419 => (x"c2",x"87",x"db",x"02"),
  1420 => (x"f7",x"c1",x"02",x"8d"),
  1421 => (x"02",x"8d",x"c9",x"87"),
  1422 => (x"c4",x"87",x"d1",x"c4"),
  1423 => (x"c2",x"c1",x"02",x"8d"),
  1424 => (x"02",x"8d",x"c1",x"87"),
  1425 => (x"c8",x"87",x"c5",x"c4"),
  1426 => (x"66",x"c8",x"87",x"e8"),
  1427 => (x"c1",x"91",x"cb",x"49"),
  1428 => (x"c4",x"81",x"66",x"c4"),
  1429 => (x"7e",x"6a",x"4a",x"a1"),
  1430 => (x"e4",x"c1",x"1e",x"71"),
  1431 => (x"66",x"c4",x"48",x"c9"),
  1432 => (x"4a",x"a1",x"cc",x"49"),
  1433 => (x"aa",x"71",x"41",x"20"),
  1434 => (x"87",x"f8",x"ff",x"05"),
  1435 => (x"49",x"26",x"51",x"10"),
  1436 => (x"79",x"f3",x"d2",x"c1"),
  1437 => (x"87",x"d5",x"dd",x"ff"),
  1438 => (x"e8",x"c0",x"4c",x"70"),
  1439 => (x"78",x"c1",x"48",x"a6"),
  1440 => (x"c4",x"87",x"f5",x"c7"),
  1441 => (x"f0",x"c0",x"48",x"a6"),
  1442 => (x"eb",x"db",x"ff",x"78"),
  1443 => (x"c0",x"4c",x"70",x"87"),
  1444 => (x"c0",x"02",x"ac",x"ec"),
  1445 => (x"a6",x"c8",x"87",x"c3"),
  1446 => (x"ac",x"ec",x"c0",x"5c"),
  1447 => (x"ff",x"87",x"cd",x"02"),
  1448 => (x"70",x"87",x"d5",x"db"),
  1449 => (x"ac",x"ec",x"c0",x"4c"),
  1450 => (x"87",x"f3",x"ff",x"05"),
  1451 => (x"02",x"ac",x"ec",x"c0"),
  1452 => (x"ff",x"87",x"c4",x"c0"),
  1453 => (x"c4",x"87",x"c1",x"db"),
  1454 => (x"66",x"d8",x"1e",x"66"),
  1455 => (x"66",x"d8",x"1e",x"49"),
  1456 => (x"e9",x"c1",x"1e",x"49"),
  1457 => (x"66",x"d8",x"1e",x"ca"),
  1458 => (x"87",x"c0",x"f8",x"49"),
  1459 => (x"1e",x"ca",x"1e",x"c0"),
  1460 => (x"49",x"66",x"e0",x"c0"),
  1461 => (x"dc",x"c1",x"91",x"cb"),
  1462 => (x"a6",x"d8",x"81",x"66"),
  1463 => (x"78",x"a1",x"c4",x"48"),
  1464 => (x"49",x"bf",x"66",x"d8"),
  1465 => (x"87",x"f9",x"db",x"ff"),
  1466 => (x"b7",x"c0",x"86",x"d8"),
  1467 => (x"cb",x"c1",x"06",x"a8"),
  1468 => (x"de",x"1e",x"c1",x"87"),
  1469 => (x"bf",x"66",x"c8",x"1e"),
  1470 => (x"e4",x"db",x"ff",x"49"),
  1471 => (x"70",x"86",x"c8",x"87"),
  1472 => (x"08",x"c0",x"48",x"49"),
  1473 => (x"a6",x"ec",x"c0",x"88"),
  1474 => (x"a8",x"b7",x"c0",x"58"),
  1475 => (x"87",x"ec",x"c0",x"06"),
  1476 => (x"48",x"66",x"e8",x"c0"),
  1477 => (x"03",x"a8",x"b7",x"dd"),
  1478 => (x"6e",x"87",x"e1",x"c0"),
  1479 => (x"e8",x"c0",x"49",x"bf"),
  1480 => (x"e0",x"c0",x"81",x"66"),
  1481 => (x"66",x"e8",x"c0",x"51"),
  1482 => (x"6e",x"81",x"c1",x"49"),
  1483 => (x"c1",x"c2",x"81",x"bf"),
  1484 => (x"66",x"e8",x"c0",x"51"),
  1485 => (x"6e",x"81",x"c2",x"49"),
  1486 => (x"51",x"c0",x"81",x"bf"),
  1487 => (x"c1",x"48",x"66",x"d0"),
  1488 => (x"58",x"a6",x"d4",x"80"),
  1489 => (x"c1",x"80",x"d8",x"48"),
  1490 => (x"87",x"ec",x"c4",x"78"),
  1491 => (x"87",x"c0",x"dc",x"ff"),
  1492 => (x"58",x"a6",x"ec",x"c0"),
  1493 => (x"87",x"f8",x"db",x"ff"),
  1494 => (x"58",x"a6",x"f0",x"c0"),
  1495 => (x"05",x"a8",x"ec",x"c0"),
  1496 => (x"a6",x"87",x"c9",x"c0"),
  1497 => (x"66",x"e8",x"c0",x"48"),
  1498 => (x"87",x"c4",x"c0",x"78"),
  1499 => (x"87",x"c8",x"d8",x"ff"),
  1500 => (x"cb",x"49",x"66",x"c8"),
  1501 => (x"66",x"c4",x"c1",x"91"),
  1502 => (x"c8",x"80",x"71",x"48"),
  1503 => (x"66",x"c4",x"58",x"a6"),
  1504 => (x"c4",x"82",x"c8",x"4a"),
  1505 => (x"81",x"ca",x"49",x"66"),
  1506 => (x"51",x"66",x"e8",x"c0"),
  1507 => (x"49",x"66",x"ec",x"c0"),
  1508 => (x"e8",x"c0",x"81",x"c1"),
  1509 => (x"48",x"c1",x"89",x"66"),
  1510 => (x"49",x"70",x"30",x"71"),
  1511 => (x"97",x"71",x"89",x"c1"),
  1512 => (x"ec",x"f8",x"c2",x"7a"),
  1513 => (x"e8",x"c0",x"49",x"bf"),
  1514 => (x"6a",x"97",x"29",x"66"),
  1515 => (x"98",x"71",x"48",x"4a"),
  1516 => (x"58",x"a6",x"f4",x"c0"),
  1517 => (x"c4",x"49",x"66",x"c4"),
  1518 => (x"c0",x"7e",x"69",x"81"),
  1519 => (x"dc",x"48",x"66",x"e0"),
  1520 => (x"c0",x"02",x"a8",x"66"),
  1521 => (x"a6",x"dc",x"87",x"c8"),
  1522 => (x"c0",x"78",x"c0",x"48"),
  1523 => (x"a6",x"dc",x"87",x"c5"),
  1524 => (x"dc",x"78",x"c1",x"48"),
  1525 => (x"e0",x"c0",x"1e",x"66"),
  1526 => (x"49",x"66",x"c8",x"1e"),
  1527 => (x"87",x"c1",x"d8",x"ff"),
  1528 => (x"4c",x"70",x"86",x"c8"),
  1529 => (x"06",x"ac",x"b7",x"c0"),
  1530 => (x"6e",x"87",x"d6",x"c1"),
  1531 => (x"70",x"80",x"74",x"48"),
  1532 => (x"49",x"e0",x"c0",x"7e"),
  1533 => (x"4b",x"6e",x"89",x"74"),
  1534 => (x"4a",x"c6",x"e4",x"c1"),
  1535 => (x"e7",x"e2",x"fe",x"71"),
  1536 => (x"c2",x"48",x"6e",x"87"),
  1537 => (x"c0",x"7e",x"70",x"80"),
  1538 => (x"c1",x"48",x"66",x"e4"),
  1539 => (x"a6",x"e8",x"c0",x"80"),
  1540 => (x"66",x"f0",x"c0",x"58"),
  1541 => (x"70",x"81",x"c1",x"49"),
  1542 => (x"c5",x"c0",x"02",x"a9"),
  1543 => (x"c0",x"4d",x"c0",x"87"),
  1544 => (x"4d",x"c1",x"87",x"c2"),
  1545 => (x"a4",x"c2",x"1e",x"75"),
  1546 => (x"48",x"e0",x"c0",x"49"),
  1547 => (x"49",x"70",x"88",x"71"),
  1548 => (x"49",x"66",x"c8",x"1e"),
  1549 => (x"87",x"e9",x"d6",x"ff"),
  1550 => (x"b7",x"c0",x"86",x"c8"),
  1551 => (x"c6",x"ff",x"01",x"a8"),
  1552 => (x"66",x"e4",x"c0",x"87"),
  1553 => (x"87",x"d3",x"c0",x"02"),
  1554 => (x"c9",x"49",x"66",x"c4"),
  1555 => (x"66",x"e4",x"c0",x"81"),
  1556 => (x"48",x"66",x"c4",x"51"),
  1557 => (x"78",x"df",x"cf",x"c1"),
  1558 => (x"c4",x"87",x"ce",x"c0"),
  1559 => (x"81",x"c9",x"49",x"66"),
  1560 => (x"66",x"c4",x"51",x"c2"),
  1561 => (x"d3",x"d0",x"c1",x"48"),
  1562 => (x"a6",x"e8",x"c0",x"78"),
  1563 => (x"c0",x"78",x"c1",x"48"),
  1564 => (x"d5",x"ff",x"87",x"c6"),
  1565 => (x"4c",x"70",x"87",x"d7"),
  1566 => (x"02",x"66",x"e8",x"c0"),
  1567 => (x"c8",x"87",x"f5",x"c0"),
  1568 => (x"66",x"cc",x"48",x"66"),
  1569 => (x"cb",x"c0",x"04",x"a8"),
  1570 => (x"48",x"66",x"c8",x"87"),
  1571 => (x"a6",x"cc",x"80",x"c1"),
  1572 => (x"87",x"e0",x"c0",x"58"),
  1573 => (x"c1",x"48",x"66",x"cc"),
  1574 => (x"58",x"a6",x"d0",x"88"),
  1575 => (x"c1",x"87",x"d5",x"c0"),
  1576 => (x"c0",x"05",x"ac",x"c6"),
  1577 => (x"66",x"d0",x"87",x"c8"),
  1578 => (x"d4",x"80",x"c1",x"48"),
  1579 => (x"d4",x"ff",x"58",x"a6"),
  1580 => (x"4c",x"70",x"87",x"db"),
  1581 => (x"c1",x"48",x"66",x"d4"),
  1582 => (x"58",x"a6",x"d8",x"80"),
  1583 => (x"c0",x"02",x"9c",x"74"),
  1584 => (x"66",x"c8",x"87",x"cb"),
  1585 => (x"66",x"cc",x"c1",x"48"),
  1586 => (x"e9",x"f3",x"04",x"a8"),
  1587 => (x"f3",x"d3",x"ff",x"87"),
  1588 => (x"48",x"66",x"c8",x"87"),
  1589 => (x"c0",x"03",x"a8",x"c7"),
  1590 => (x"f5",x"c2",x"87",x"e5"),
  1591 => (x"78",x"c0",x"48",x"c0"),
  1592 => (x"cb",x"49",x"66",x"c8"),
  1593 => (x"66",x"c4",x"c1",x"91"),
  1594 => (x"4a",x"a1",x"c4",x"81"),
  1595 => (x"52",x"c0",x"4a",x"6a"),
  1596 => (x"48",x"66",x"c8",x"79"),
  1597 => (x"a6",x"cc",x"80",x"c1"),
  1598 => (x"04",x"a8",x"c7",x"58"),
  1599 => (x"ff",x"87",x"db",x"ff"),
  1600 => (x"df",x"ff",x"8e",x"cc"),
  1601 => (x"20",x"3a",x"87",x"f7"),
  1602 => (x"50",x"49",x"44",x"00"),
  1603 => (x"69",x"77",x"53",x"20"),
  1604 => (x"65",x"68",x"63",x"74"),
  1605 => (x"73",x"1e",x"00",x"73"),
  1606 => (x"9b",x"4b",x"71",x"1e"),
  1607 => (x"c2",x"87",x"c6",x"02"),
  1608 => (x"c0",x"48",x"fc",x"f4"),
  1609 => (x"c2",x"1e",x"c7",x"78"),
  1610 => (x"49",x"bf",x"fc",x"f4"),
  1611 => (x"e7",x"e7",x"c1",x"1e"),
  1612 => (x"e4",x"f4",x"c2",x"1e"),
  1613 => (x"c8",x"ef",x"49",x"bf"),
  1614 => (x"c2",x"86",x"cc",x"87"),
  1615 => (x"49",x"bf",x"e4",x"f4"),
  1616 => (x"73",x"87",x"f4",x"e9"),
  1617 => (x"87",x"c8",x"02",x"9b"),
  1618 => (x"49",x"e7",x"e7",x"c1"),
  1619 => (x"87",x"f7",x"ed",x"c0"),
  1620 => (x"87",x"ed",x"de",x"ff"),
  1621 => (x"87",x"d1",x"c7",x"1e"),
  1622 => (x"f9",x"fe",x"49",x"c1"),
  1623 => (x"e2",x"e5",x"fe",x"87"),
  1624 => (x"02",x"98",x"70",x"87"),
  1625 => (x"ec",x"fe",x"87",x"cd"),
  1626 => (x"98",x"70",x"87",x"fb"),
  1627 => (x"c1",x"87",x"c4",x"02"),
  1628 => (x"c0",x"87",x"c2",x"4a"),
  1629 => (x"05",x"9a",x"72",x"4a"),
  1630 => (x"1e",x"c0",x"87",x"ce"),
  1631 => (x"49",x"e9",x"e6",x"c1"),
  1632 => (x"87",x"e1",x"f9",x"c0"),
  1633 => (x"87",x"fe",x"86",x"c4"),
  1634 => (x"87",x"c4",x"fc",x"c0"),
  1635 => (x"e6",x"c1",x"1e",x"c0"),
  1636 => (x"f9",x"c0",x"49",x"f4"),
  1637 => (x"1e",x"c0",x"87",x"cf"),
  1638 => (x"87",x"ca",x"fe",x"c0"),
  1639 => (x"f9",x"c0",x"49",x"70"),
  1640 => (x"c3",x"c3",x"87",x"c3"),
  1641 => (x"26",x"8e",x"f8",x"87"),
  1642 => (x"20",x"44",x"53",x"4f"),
  1643 => (x"6c",x"69",x"61",x"66"),
  1644 => (x"00",x"2e",x"64",x"65"),
  1645 => (x"74",x"6f",x"6f",x"42"),
  1646 => (x"2e",x"67",x"6e",x"69"),
  1647 => (x"1e",x"00",x"2e",x"2e"),
  1648 => (x"48",x"fc",x"f4",x"c2"),
  1649 => (x"f4",x"c2",x"78",x"c0"),
  1650 => (x"78",x"c0",x"48",x"e4"),
  1651 => (x"c0",x"87",x"c5",x"fe"),
  1652 => (x"c0",x"87",x"e5",x"ff"),
  1653 => (x"00",x"4f",x"26",x"48"),
  1654 => (x"45",x"20",x"80",x"00"),
  1655 => (x"00",x"74",x"69",x"78"),
  1656 => (x"61",x"42",x"20",x"80"),
  1657 => (x"8f",x"00",x"6b",x"63"),
  1658 => (x"50",x"00",x"00",x"13"),
  1659 => (x"00",x"00",x"00",x"2d"),
  1660 => (x"13",x"8f",x"00",x"00"),
  1661 => (x"2d",x"6e",x"00",x"00"),
  1662 => (x"00",x"00",x"00",x"00"),
  1663 => (x"00",x"13",x"8f",x"00"),
  1664 => (x"00",x"2d",x"8c",x"00"),
  1665 => (x"00",x"00",x"00",x"00"),
  1666 => (x"00",x"00",x"13",x"8f"),
  1667 => (x"00",x"00",x"2d",x"aa"),
  1668 => (x"8f",x"00",x"00",x"00"),
  1669 => (x"c8",x"00",x"00",x"13"),
  1670 => (x"00",x"00",x"00",x"2d"),
  1671 => (x"13",x"8f",x"00",x"00"),
  1672 => (x"2d",x"e6",x"00",x"00"),
  1673 => (x"00",x"00",x"00",x"00"),
  1674 => (x"00",x"13",x"8f",x"00"),
  1675 => (x"00",x"2e",x"04",x"00"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"00",x"00",x"13",x"8f"),
  1678 => (x"00",x"00",x"00",x"00"),
  1679 => (x"24",x"00",x"00",x"00"),
  1680 => (x"00",x"00",x"00",x"14"),
  1681 => (x"00",x"00",x"00",x"00"),
  1682 => (x"6f",x"4c",x"00",x"00"),
  1683 => (x"2a",x"20",x"64",x"61"),
  1684 => (x"fe",x"1e",x"00",x"2e"),
  1685 => (x"78",x"c0",x"48",x"f0"),
  1686 => (x"09",x"79",x"09",x"cd"),
  1687 => (x"1e",x"1e",x"4f",x"26"),
  1688 => (x"7e",x"bf",x"f0",x"fe"),
  1689 => (x"4f",x"26",x"26",x"48"),
  1690 => (x"48",x"f0",x"fe",x"1e"),
  1691 => (x"4f",x"26",x"78",x"c1"),
  1692 => (x"48",x"f0",x"fe",x"1e"),
  1693 => (x"4f",x"26",x"78",x"c0"),
  1694 => (x"c0",x"4a",x"71",x"1e"),
  1695 => (x"4f",x"26",x"52",x"52"),
  1696 => (x"5c",x"5b",x"5e",x"0e"),
  1697 => (x"86",x"f4",x"0e",x"5d"),
  1698 => (x"6d",x"97",x"4d",x"71"),
  1699 => (x"4c",x"a5",x"c1",x"7e"),
  1700 => (x"c8",x"48",x"6c",x"97"),
  1701 => (x"48",x"6e",x"58",x"a6"),
  1702 => (x"05",x"a8",x"66",x"c4"),
  1703 => (x"48",x"ff",x"87",x"c5"),
  1704 => (x"ff",x"87",x"e6",x"c0"),
  1705 => (x"a5",x"c2",x"87",x"ca"),
  1706 => (x"4b",x"6c",x"97",x"49"),
  1707 => (x"97",x"4b",x"a3",x"71"),
  1708 => (x"6c",x"97",x"4b",x"6b"),
  1709 => (x"c1",x"48",x"6e",x"7e"),
  1710 => (x"58",x"a6",x"c8",x"80"),
  1711 => (x"a6",x"cc",x"98",x"c7"),
  1712 => (x"7c",x"97",x"70",x"58"),
  1713 => (x"73",x"87",x"e1",x"fe"),
  1714 => (x"26",x"8e",x"f4",x"48"),
  1715 => (x"26",x"4c",x"26",x"4d"),
  1716 => (x"0e",x"4f",x"26",x"4b"),
  1717 => (x"0e",x"5c",x"5b",x"5e"),
  1718 => (x"4c",x"71",x"86",x"f4"),
  1719 => (x"c3",x"4a",x"66",x"d8"),
  1720 => (x"a4",x"c2",x"9a",x"ff"),
  1721 => (x"49",x"6c",x"97",x"4b"),
  1722 => (x"72",x"49",x"a1",x"73"),
  1723 => (x"7e",x"6c",x"97",x"51"),
  1724 => (x"80",x"c1",x"48",x"6e"),
  1725 => (x"c7",x"58",x"a6",x"c8"),
  1726 => (x"58",x"a6",x"cc",x"98"),
  1727 => (x"8e",x"f4",x"54",x"70"),
  1728 => (x"1e",x"87",x"ca",x"ff"),
  1729 => (x"87",x"e8",x"fd",x"1e"),
  1730 => (x"49",x"4a",x"bf",x"e0"),
  1731 => (x"99",x"c0",x"e0",x"c0"),
  1732 => (x"72",x"87",x"cb",x"02"),
  1733 => (x"e2",x"f8",x"c2",x"1e"),
  1734 => (x"87",x"f7",x"fe",x"49"),
  1735 => (x"fd",x"fc",x"86",x"c4"),
  1736 => (x"fd",x"7e",x"70",x"87"),
  1737 => (x"26",x"26",x"87",x"c2"),
  1738 => (x"f8",x"c2",x"1e",x"4f"),
  1739 => (x"c7",x"fd",x"49",x"e2"),
  1740 => (x"c3",x"ec",x"c1",x"87"),
  1741 => (x"87",x"da",x"fc",x"49"),
  1742 => (x"26",x"87",x"c8",x"c4"),
  1743 => (x"d0",x"ff",x"1e",x"4f"),
  1744 => (x"78",x"e1",x"c8",x"48"),
  1745 => (x"c5",x"48",x"d4",x"ff"),
  1746 => (x"02",x"66",x"c4",x"78"),
  1747 => (x"e0",x"c3",x"87",x"c3"),
  1748 => (x"02",x"66",x"c8",x"78"),
  1749 => (x"d4",x"ff",x"87",x"c6"),
  1750 => (x"78",x"f0",x"c3",x"48"),
  1751 => (x"71",x"48",x"d4",x"ff"),
  1752 => (x"48",x"d0",x"ff",x"78"),
  1753 => (x"c0",x"78",x"e1",x"c8"),
  1754 => (x"4f",x"26",x"78",x"e0"),
  1755 => (x"5c",x"5b",x"5e",x"0e"),
  1756 => (x"c2",x"4c",x"71",x"0e"),
  1757 => (x"fc",x"49",x"e2",x"f8"),
  1758 => (x"4a",x"70",x"87",x"c6"),
  1759 => (x"04",x"aa",x"b7",x"c0"),
  1760 => (x"c3",x"87",x"e3",x"c2"),
  1761 => (x"c9",x"05",x"aa",x"e0"),
  1762 => (x"f6",x"f0",x"c1",x"87"),
  1763 => (x"c2",x"78",x"c1",x"48"),
  1764 => (x"f0",x"c3",x"87",x"d4"),
  1765 => (x"87",x"c9",x"05",x"aa"),
  1766 => (x"48",x"f2",x"f0",x"c1"),
  1767 => (x"f5",x"c1",x"78",x"c1"),
  1768 => (x"f6",x"f0",x"c1",x"87"),
  1769 => (x"87",x"c7",x"02",x"bf"),
  1770 => (x"c0",x"c2",x"4b",x"72"),
  1771 => (x"72",x"87",x"c2",x"b3"),
  1772 => (x"05",x"9c",x"74",x"4b"),
  1773 => (x"f0",x"c1",x"87",x"d1"),
  1774 => (x"c1",x"1e",x"bf",x"f2"),
  1775 => (x"1e",x"bf",x"f6",x"f0"),
  1776 => (x"f8",x"fd",x"49",x"72"),
  1777 => (x"c1",x"86",x"c8",x"87"),
  1778 => (x"02",x"bf",x"f2",x"f0"),
  1779 => (x"73",x"87",x"e0",x"c0"),
  1780 => (x"29",x"b7",x"c4",x"49"),
  1781 => (x"d2",x"f2",x"c1",x"91"),
  1782 => (x"cf",x"4a",x"73",x"81"),
  1783 => (x"c1",x"92",x"c2",x"9a"),
  1784 => (x"70",x"30",x"72",x"48"),
  1785 => (x"72",x"ba",x"ff",x"4a"),
  1786 => (x"70",x"98",x"69",x"48"),
  1787 => (x"73",x"87",x"db",x"79"),
  1788 => (x"29",x"b7",x"c4",x"49"),
  1789 => (x"d2",x"f2",x"c1",x"91"),
  1790 => (x"cf",x"4a",x"73",x"81"),
  1791 => (x"c3",x"92",x"c2",x"9a"),
  1792 => (x"70",x"30",x"72",x"48"),
  1793 => (x"b0",x"69",x"48",x"4a"),
  1794 => (x"f0",x"c1",x"79",x"70"),
  1795 => (x"78",x"c0",x"48",x"f6"),
  1796 => (x"48",x"f2",x"f0",x"c1"),
  1797 => (x"f8",x"c2",x"78",x"c0"),
  1798 => (x"e3",x"f9",x"49",x"e2"),
  1799 => (x"c0",x"4a",x"70",x"87"),
  1800 => (x"fd",x"03",x"aa",x"b7"),
  1801 => (x"48",x"c0",x"87",x"dd"),
  1802 => (x"4d",x"26",x"87",x"c2"),
  1803 => (x"4b",x"26",x"4c",x"26"),
  1804 => (x"00",x"00",x"4f",x"26"),
  1805 => (x"00",x"00",x"00",x"00"),
  1806 => (x"71",x"1e",x"00",x"00"),
  1807 => (x"eb",x"fc",x"49",x"4a"),
  1808 => (x"1e",x"4f",x"26",x"87"),
  1809 => (x"49",x"72",x"4a",x"c0"),
  1810 => (x"f2",x"c1",x"91",x"c4"),
  1811 => (x"79",x"c0",x"81",x"d2"),
  1812 => (x"b7",x"d0",x"82",x"c1"),
  1813 => (x"87",x"ee",x"04",x"aa"),
  1814 => (x"5e",x"0e",x"4f",x"26"),
  1815 => (x"0e",x"5d",x"5c",x"5b"),
  1816 => (x"cb",x"f8",x"4d",x"71"),
  1817 => (x"c4",x"4a",x"75",x"87"),
  1818 => (x"c1",x"92",x"2a",x"b7"),
  1819 => (x"75",x"82",x"d2",x"f2"),
  1820 => (x"c2",x"9c",x"cf",x"4c"),
  1821 => (x"4b",x"49",x"6a",x"94"),
  1822 => (x"9b",x"c3",x"2b",x"74"),
  1823 => (x"30",x"74",x"48",x"c2"),
  1824 => (x"bc",x"ff",x"4c",x"70"),
  1825 => (x"98",x"71",x"48",x"74"),
  1826 => (x"db",x"f7",x"7a",x"70"),
  1827 => (x"fe",x"48",x"73",x"87"),
  1828 => (x"00",x"00",x"87",x"d8"),
  1829 => (x"00",x"00",x"00",x"00"),
  1830 => (x"00",x"00",x"00",x"00"),
  1831 => (x"00",x"00",x"00",x"00"),
  1832 => (x"00",x"00",x"00",x"00"),
  1833 => (x"00",x"00",x"00",x"00"),
  1834 => (x"00",x"00",x"00",x"00"),
  1835 => (x"00",x"00",x"00",x"00"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"00",x"00",x"00",x"00"),
  1838 => (x"00",x"00",x"00",x"00"),
  1839 => (x"00",x"00",x"00",x"00"),
  1840 => (x"00",x"00",x"00",x"00"),
  1841 => (x"00",x"00",x"00",x"00"),
  1842 => (x"00",x"00",x"00",x"00"),
  1843 => (x"00",x"00",x"00",x"00"),
  1844 => (x"ff",x"1e",x"00",x"00"),
  1845 => (x"e1",x"c8",x"48",x"d0"),
  1846 => (x"ff",x"48",x"71",x"78"),
  1847 => (x"c4",x"78",x"08",x"d4"),
  1848 => (x"d4",x"ff",x"48",x"66"),
  1849 => (x"4f",x"26",x"78",x"08"),
  1850 => (x"c4",x"4a",x"71",x"1e"),
  1851 => (x"72",x"1e",x"49",x"66"),
  1852 => (x"87",x"de",x"ff",x"49"),
  1853 => (x"c0",x"48",x"d0",x"ff"),
  1854 => (x"26",x"26",x"78",x"e0"),
  1855 => (x"1e",x"73",x"1e",x"4f"),
  1856 => (x"66",x"c8",x"4b",x"71"),
  1857 => (x"4a",x"73",x"1e",x"49"),
  1858 => (x"49",x"a2",x"e0",x"c1"),
  1859 => (x"26",x"87",x"d9",x"ff"),
  1860 => (x"4d",x"26",x"87",x"c4"),
  1861 => (x"4b",x"26",x"4c",x"26"),
  1862 => (x"ff",x"1e",x"4f",x"26"),
  1863 => (x"ff",x"c3",x"4a",x"d4"),
  1864 => (x"48",x"d0",x"ff",x"7a"),
  1865 => (x"de",x"78",x"e1",x"c0"),
  1866 => (x"ec",x"f8",x"c2",x"7a"),
  1867 => (x"48",x"49",x"7a",x"bf"),
  1868 => (x"7a",x"70",x"28",x"c8"),
  1869 => (x"28",x"d0",x"48",x"71"),
  1870 => (x"48",x"71",x"7a",x"70"),
  1871 => (x"7a",x"70",x"28",x"d8"),
  1872 => (x"c0",x"48",x"d0",x"ff"),
  1873 => (x"4f",x"26",x"78",x"e0"),
  1874 => (x"5c",x"5b",x"5e",x"0e"),
  1875 => (x"4c",x"71",x"0e",x"5d"),
  1876 => (x"bf",x"ec",x"f8",x"c2"),
  1877 => (x"2b",x"74",x"4b",x"4d"),
  1878 => (x"c1",x"9b",x"66",x"d0"),
  1879 => (x"ab",x"66",x"d4",x"83"),
  1880 => (x"c0",x"87",x"c2",x"04"),
  1881 => (x"d0",x"4a",x"74",x"4b"),
  1882 => (x"31",x"72",x"49",x"66"),
  1883 => (x"99",x"75",x"b9",x"ff"),
  1884 => (x"30",x"72",x"48",x"73"),
  1885 => (x"71",x"48",x"4a",x"70"),
  1886 => (x"f0",x"f8",x"c2",x"b0"),
  1887 => (x"87",x"da",x"fe",x"58"),
  1888 => (x"4c",x"26",x"4d",x"26"),
  1889 => (x"4f",x"26",x"4b",x"26"),
  1890 => (x"5c",x"5b",x"5e",x"0e"),
  1891 => (x"71",x"1e",x"0e",x"5d"),
  1892 => (x"f0",x"f8",x"c2",x"4c"),
  1893 => (x"c0",x"4a",x"c0",x"4b"),
  1894 => (x"cc",x"fe",x"49",x"f4"),
  1895 => (x"1e",x"74",x"87",x"e7"),
  1896 => (x"49",x"f0",x"f8",x"c2"),
  1897 => (x"87",x"c9",x"e9",x"fe"),
  1898 => (x"49",x"70",x"86",x"c4"),
  1899 => (x"ea",x"c0",x"02",x"99"),
  1900 => (x"a6",x"1e",x"c4",x"87"),
  1901 => (x"f8",x"c2",x"1e",x"4d"),
  1902 => (x"ee",x"fe",x"49",x"f0"),
  1903 => (x"86",x"c8",x"87",x"fe"),
  1904 => (x"d6",x"02",x"98",x"70"),
  1905 => (x"c1",x"4a",x"75",x"87"),
  1906 => (x"c4",x"49",x"d1",x"f8"),
  1907 => (x"d9",x"ca",x"fe",x"4b"),
  1908 => (x"02",x"98",x"70",x"87"),
  1909 => (x"48",x"c0",x"87",x"ca"),
  1910 => (x"c0",x"87",x"ed",x"c0"),
  1911 => (x"87",x"e8",x"c0",x"48"),
  1912 => (x"c1",x"87",x"f3",x"c0"),
  1913 => (x"98",x"70",x"87",x"c4"),
  1914 => (x"c0",x"87",x"c8",x"02"),
  1915 => (x"98",x"70",x"87",x"fc"),
  1916 => (x"c2",x"87",x"f8",x"05"),
  1917 => (x"02",x"bf",x"d0",x"f9"),
  1918 => (x"f8",x"c2",x"87",x"cc"),
  1919 => (x"f9",x"c2",x"48",x"ec"),
  1920 => (x"fc",x"78",x"bf",x"d0"),
  1921 => (x"48",x"c1",x"87",x"d4"),
  1922 => (x"26",x"4d",x"26",x"26"),
  1923 => (x"26",x"4b",x"26",x"4c"),
  1924 => (x"52",x"41",x"5b",x"4f"),
  1925 => (x"c0",x"1e",x"00",x"43"),
  1926 => (x"f0",x"f8",x"c2",x"1e"),
  1927 => (x"f4",x"eb",x"fe",x"49"),
  1928 => (x"c8",x"f9",x"c2",x"87"),
  1929 => (x"26",x"78",x"c0",x"48"),
  1930 => (x"5e",x"0e",x"4f",x"26"),
  1931 => (x"0e",x"5d",x"5c",x"5b"),
  1932 => (x"a6",x"c4",x"86",x"f4"),
  1933 => (x"c2",x"78",x"c0",x"48"),
  1934 => (x"48",x"bf",x"c8",x"f9"),
  1935 => (x"03",x"a8",x"b7",x"c3"),
  1936 => (x"f9",x"c2",x"87",x"d1"),
  1937 => (x"c1",x"48",x"bf",x"c8"),
  1938 => (x"cc",x"f9",x"c2",x"80"),
  1939 => (x"48",x"fb",x"c0",x"58"),
  1940 => (x"c2",x"87",x"e2",x"c6"),
  1941 => (x"fe",x"49",x"f0",x"f8"),
  1942 => (x"70",x"87",x"f5",x"f0"),
  1943 => (x"c8",x"f9",x"c2",x"4c"),
  1944 => (x"8a",x"c3",x"4a",x"bf"),
  1945 => (x"c1",x"87",x"d8",x"02"),
  1946 => (x"cb",x"c5",x"02",x"8a"),
  1947 => (x"c2",x"02",x"8a",x"87"),
  1948 => (x"02",x"8a",x"87",x"f6"),
  1949 => (x"8a",x"87",x"cd",x"c1"),
  1950 => (x"87",x"e2",x"c3",x"02"),
  1951 => (x"c0",x"87",x"e1",x"c5"),
  1952 => (x"c4",x"4a",x"75",x"4d"),
  1953 => (x"d3",x"c0",x"c2",x"92"),
  1954 => (x"c4",x"f9",x"c2",x"82"),
  1955 => (x"70",x"80",x"75",x"48"),
  1956 => (x"bf",x"97",x"6e",x"7e"),
  1957 => (x"6e",x"4b",x"49",x"4b"),
  1958 => (x"50",x"a3",x"c1",x"48"),
  1959 => (x"48",x"11",x"81",x"6a"),
  1960 => (x"70",x"58",x"a6",x"cc"),
  1961 => (x"87",x"c4",x"02",x"ac"),
  1962 => (x"50",x"c0",x"48",x"6e"),
  1963 => (x"c7",x"05",x"66",x"c8"),
  1964 => (x"c8",x"f9",x"c2",x"87"),
  1965 => (x"78",x"a5",x"c4",x"48"),
  1966 => (x"b7",x"c4",x"85",x"c1"),
  1967 => (x"c0",x"ff",x"04",x"ad"),
  1968 => (x"87",x"dc",x"c4",x"87"),
  1969 => (x"bf",x"d4",x"f9",x"c2"),
  1970 => (x"a8",x"b7",x"c8",x"48"),
  1971 => (x"ca",x"87",x"d1",x"01"),
  1972 => (x"87",x"cc",x"02",x"ac"),
  1973 => (x"c7",x"02",x"ac",x"cd"),
  1974 => (x"ac",x"b7",x"c0",x"87"),
  1975 => (x"87",x"f3",x"c0",x"03"),
  1976 => (x"bf",x"d4",x"f9",x"c2"),
  1977 => (x"ab",x"b7",x"c8",x"4b"),
  1978 => (x"c2",x"87",x"d2",x"03"),
  1979 => (x"73",x"49",x"d8",x"f9"),
  1980 => (x"51",x"e0",x"c0",x"81"),
  1981 => (x"b7",x"c8",x"83",x"c1"),
  1982 => (x"ee",x"ff",x"04",x"ab"),
  1983 => (x"e0",x"f9",x"c2",x"87"),
  1984 => (x"50",x"d2",x"c1",x"48"),
  1985 => (x"c1",x"50",x"cf",x"c1"),
  1986 => (x"50",x"c0",x"50",x"cd"),
  1987 => (x"78",x"c3",x"80",x"e4"),
  1988 => (x"c2",x"87",x"cd",x"c3"),
  1989 => (x"49",x"bf",x"d4",x"f9"),
  1990 => (x"c2",x"80",x"c1",x"48"),
  1991 => (x"48",x"58",x"d8",x"f9"),
  1992 => (x"74",x"81",x"a0",x"c4"),
  1993 => (x"87",x"f8",x"c2",x"51"),
  1994 => (x"ac",x"b7",x"f0",x"c0"),
  1995 => (x"c0",x"87",x"da",x"04"),
  1996 => (x"01",x"ac",x"b7",x"f9"),
  1997 => (x"f9",x"c2",x"87",x"d3"),
  1998 => (x"ca",x"49",x"bf",x"cc"),
  1999 => (x"c0",x"4a",x"74",x"91"),
  2000 => (x"f9",x"c2",x"8a",x"f0"),
  2001 => (x"a1",x"72",x"48",x"cc"),
  2002 => (x"02",x"ac",x"ca",x"78"),
  2003 => (x"cd",x"87",x"c6",x"c0"),
  2004 => (x"cb",x"c2",x"05",x"ac"),
  2005 => (x"c8",x"f9",x"c2",x"87"),
  2006 => (x"c2",x"78",x"c3",x"48"),
  2007 => (x"f0",x"c0",x"87",x"c2"),
  2008 => (x"db",x"04",x"ac",x"b7"),
  2009 => (x"b7",x"f9",x"c0",x"87"),
  2010 => (x"d3",x"c0",x"01",x"ac"),
  2011 => (x"d0",x"f9",x"c2",x"87"),
  2012 => (x"91",x"d0",x"49",x"bf"),
  2013 => (x"f0",x"c0",x"4a",x"74"),
  2014 => (x"d0",x"f9",x"c2",x"8a"),
  2015 => (x"78",x"a1",x"72",x"48"),
  2016 => (x"ac",x"b7",x"c1",x"c1"),
  2017 => (x"87",x"db",x"c0",x"04"),
  2018 => (x"ac",x"b7",x"c6",x"c1"),
  2019 => (x"87",x"d3",x"c0",x"01"),
  2020 => (x"bf",x"d0",x"f9",x"c2"),
  2021 => (x"74",x"91",x"d0",x"49"),
  2022 => (x"8a",x"f7",x"c0",x"4a"),
  2023 => (x"48",x"d0",x"f9",x"c2"),
  2024 => (x"ca",x"78",x"a1",x"72"),
  2025 => (x"c6",x"c0",x"02",x"ac"),
  2026 => (x"05",x"ac",x"cd",x"87"),
  2027 => (x"c2",x"87",x"f1",x"c0"),
  2028 => (x"c3",x"48",x"c8",x"f9"),
  2029 => (x"87",x"e8",x"c0",x"78"),
  2030 => (x"05",x"ac",x"e2",x"c0"),
  2031 => (x"c4",x"87",x"c9",x"c0"),
  2032 => (x"fb",x"c0",x"48",x"a6"),
  2033 => (x"87",x"d8",x"c0",x"78"),
  2034 => (x"c0",x"02",x"ac",x"ca"),
  2035 => (x"ac",x"cd",x"87",x"c6"),
  2036 => (x"87",x"c9",x"c0",x"05"),
  2037 => (x"48",x"c8",x"f9",x"c2"),
  2038 => (x"c3",x"c0",x"78",x"c3"),
  2039 => (x"5c",x"a6",x"c8",x"87"),
  2040 => (x"03",x"ac",x"b7",x"c0"),
  2041 => (x"48",x"87",x"c4",x"c0"),
  2042 => (x"c4",x"87",x"ca",x"c0"),
  2043 => (x"c6",x"f9",x"02",x"66"),
  2044 => (x"ff",x"c3",x"48",x"87"),
  2045 => (x"f8",x"8e",x"f4",x"99"),
  2046 => (x"4f",x"43",x"87",x"cf"),
  2047 => (x"00",x"3d",x"46",x"4e"),
  2048 => (x"00",x"44",x"4f",x"4d"),
  2049 => (x"45",x"4d",x"41",x"4e"),
  2050 => (x"46",x"45",x"44",x"00"),
  2051 => (x"54",x"4c",x"55",x"41"),
  2052 => (x"fa",x"00",x"30",x"3d"),
  2053 => (x"00",x"00",x"00",x"1f"),
  2054 => (x"04",x"00",x"00",x"20"),
  2055 => (x"09",x"00",x"00",x"20"),
  2056 => (x"1e",x"00",x"00",x"20"),
  2057 => (x"c8",x"48",x"d0",x"ff"),
  2058 => (x"48",x"71",x"78",x"c9"),
  2059 => (x"78",x"08",x"d4",x"ff"),
  2060 => (x"71",x"1e",x"4f",x"26"),
  2061 => (x"87",x"eb",x"49",x"4a"),
  2062 => (x"c8",x"48",x"d0",x"ff"),
  2063 => (x"1e",x"4f",x"26",x"78"),
  2064 => (x"4b",x"71",x"1e",x"73"),
  2065 => (x"bf",x"f0",x"f9",x"c2"),
  2066 => (x"c2",x"87",x"c3",x"02"),
  2067 => (x"d0",x"ff",x"87",x"eb"),
  2068 => (x"78",x"c9",x"c8",x"48"),
  2069 => (x"e0",x"c0",x"49",x"73"),
  2070 => (x"48",x"d4",x"ff",x"b1"),
  2071 => (x"f9",x"c2",x"78",x"71"),
  2072 => (x"78",x"c0",x"48",x"e4"),
  2073 => (x"c5",x"02",x"66",x"c8"),
  2074 => (x"49",x"ff",x"c3",x"87"),
  2075 => (x"49",x"c0",x"87",x"c2"),
  2076 => (x"59",x"ec",x"f9",x"c2"),
  2077 => (x"c6",x"02",x"66",x"cc"),
  2078 => (x"d5",x"d5",x"c5",x"87"),
  2079 => (x"cf",x"87",x"c4",x"4a"),
  2080 => (x"c2",x"4a",x"ff",x"ff"),
  2081 => (x"c2",x"5a",x"f0",x"f9"),
  2082 => (x"c1",x"48",x"f0",x"f9"),
  2083 => (x"26",x"87",x"c4",x"78"),
  2084 => (x"26",x"4c",x"26",x"4d"),
  2085 => (x"0e",x"4f",x"26",x"4b"),
  2086 => (x"5d",x"5c",x"5b",x"5e"),
  2087 => (x"c2",x"4a",x"71",x"0e"),
  2088 => (x"4c",x"bf",x"ec",x"f9"),
  2089 => (x"cb",x"02",x"9a",x"72"),
  2090 => (x"91",x"c8",x"49",x"87"),
  2091 => (x"4b",x"f5",x"c0",x"c2"),
  2092 => (x"87",x"c4",x"83",x"71"),
  2093 => (x"4b",x"f5",x"c4",x"c2"),
  2094 => (x"49",x"13",x"4d",x"c0"),
  2095 => (x"f9",x"c2",x"99",x"74"),
  2096 => (x"ff",x"b9",x"bf",x"e8"),
  2097 => (x"78",x"71",x"48",x"d4"),
  2098 => (x"85",x"2c",x"b7",x"c1"),
  2099 => (x"04",x"ad",x"b7",x"c8"),
  2100 => (x"f9",x"c2",x"87",x"e8"),
  2101 => (x"c8",x"48",x"bf",x"e4"),
  2102 => (x"e8",x"f9",x"c2",x"80"),
  2103 => (x"87",x"ef",x"fe",x"58"),
  2104 => (x"71",x"1e",x"73",x"1e"),
  2105 => (x"9a",x"4a",x"13",x"4b"),
  2106 => (x"72",x"87",x"cb",x"02"),
  2107 => (x"87",x"e7",x"fe",x"49"),
  2108 => (x"05",x"9a",x"4a",x"13"),
  2109 => (x"da",x"fe",x"87",x"f5"),
  2110 => (x"f9",x"c2",x"1e",x"87"),
  2111 => (x"c2",x"49",x"bf",x"e4"),
  2112 => (x"c1",x"48",x"e4",x"f9"),
  2113 => (x"c0",x"c4",x"78",x"a1"),
  2114 => (x"db",x"03",x"a9",x"b7"),
  2115 => (x"48",x"d4",x"ff",x"87"),
  2116 => (x"bf",x"e8",x"f9",x"c2"),
  2117 => (x"e4",x"f9",x"c2",x"78"),
  2118 => (x"f9",x"c2",x"49",x"bf"),
  2119 => (x"a1",x"c1",x"48",x"e4"),
  2120 => (x"b7",x"c0",x"c4",x"78"),
  2121 => (x"87",x"e5",x"04",x"a9"),
  2122 => (x"c8",x"48",x"d0",x"ff"),
  2123 => (x"f0",x"f9",x"c2",x"78"),
  2124 => (x"26",x"78",x"c0",x"48"),
  2125 => (x"00",x"00",x"00",x"4f"),
  2126 => (x"00",x"00",x"00",x"00"),
  2127 => (x"00",x"00",x"00",x"00"),
  2128 => (x"00",x"00",x"5f",x"5f"),
  2129 => (x"03",x"03",x"00",x"00"),
  2130 => (x"00",x"03",x"03",x"00"),
  2131 => (x"7f",x"7f",x"14",x"00"),
  2132 => (x"14",x"7f",x"7f",x"14"),
  2133 => (x"2e",x"24",x"00",x"00"),
  2134 => (x"12",x"3a",x"6b",x"6b"),
  2135 => (x"36",x"6a",x"4c",x"00"),
  2136 => (x"32",x"56",x"6c",x"18"),
  2137 => (x"4f",x"7e",x"30",x"00"),
  2138 => (x"68",x"3a",x"77",x"59"),
  2139 => (x"04",x"00",x"00",x"40"),
  2140 => (x"00",x"00",x"03",x"07"),
  2141 => (x"1c",x"00",x"00",x"00"),
  2142 => (x"00",x"41",x"63",x"3e"),
  2143 => (x"41",x"00",x"00",x"00"),
  2144 => (x"00",x"1c",x"3e",x"63"),
  2145 => (x"3e",x"2a",x"08",x"00"),
  2146 => (x"2a",x"3e",x"1c",x"1c"),
  2147 => (x"08",x"08",x"00",x"08"),
  2148 => (x"08",x"08",x"3e",x"3e"),
  2149 => (x"80",x"00",x"00",x"00"),
  2150 => (x"00",x"00",x"60",x"e0"),
  2151 => (x"08",x"08",x"00",x"00"),
  2152 => (x"08",x"08",x"08",x"08"),
  2153 => (x"00",x"00",x"00",x"00"),
  2154 => (x"00",x"00",x"60",x"60"),
  2155 => (x"30",x"60",x"40",x"00"),
  2156 => (x"03",x"06",x"0c",x"18"),
  2157 => (x"7f",x"3e",x"00",x"01"),
  2158 => (x"3e",x"7f",x"4d",x"59"),
  2159 => (x"06",x"04",x"00",x"00"),
  2160 => (x"00",x"00",x"7f",x"7f"),
  2161 => (x"63",x"42",x"00",x"00"),
  2162 => (x"46",x"4f",x"59",x"71"),
  2163 => (x"63",x"22",x"00",x"00"),
  2164 => (x"36",x"7f",x"49",x"49"),
  2165 => (x"16",x"1c",x"18",x"00"),
  2166 => (x"10",x"7f",x"7f",x"13"),
  2167 => (x"67",x"27",x"00",x"00"),
  2168 => (x"39",x"7d",x"45",x"45"),
  2169 => (x"7e",x"3c",x"00",x"00"),
  2170 => (x"30",x"79",x"49",x"4b"),
  2171 => (x"01",x"01",x"00",x"00"),
  2172 => (x"07",x"0f",x"79",x"71"),
  2173 => (x"7f",x"36",x"00",x"00"),
  2174 => (x"36",x"7f",x"49",x"49"),
  2175 => (x"4f",x"06",x"00",x"00"),
  2176 => (x"1e",x"3f",x"69",x"49"),
  2177 => (x"00",x"00",x"00",x"00"),
  2178 => (x"00",x"00",x"66",x"66"),
  2179 => (x"80",x"00",x"00",x"00"),
  2180 => (x"00",x"00",x"66",x"e6"),
  2181 => (x"08",x"08",x"00",x"00"),
  2182 => (x"22",x"22",x"14",x"14"),
  2183 => (x"14",x"14",x"00",x"00"),
  2184 => (x"14",x"14",x"14",x"14"),
  2185 => (x"22",x"22",x"00",x"00"),
  2186 => (x"08",x"08",x"14",x"14"),
  2187 => (x"03",x"02",x"00",x"00"),
  2188 => (x"06",x"0f",x"59",x"51"),
  2189 => (x"41",x"7f",x"3e",x"00"),
  2190 => (x"1e",x"1f",x"55",x"5d"),
  2191 => (x"7f",x"7e",x"00",x"00"),
  2192 => (x"7e",x"7f",x"09",x"09"),
  2193 => (x"7f",x"7f",x"00",x"00"),
  2194 => (x"36",x"7f",x"49",x"49"),
  2195 => (x"3e",x"1c",x"00",x"00"),
  2196 => (x"41",x"41",x"41",x"63"),
  2197 => (x"7f",x"7f",x"00",x"00"),
  2198 => (x"1c",x"3e",x"63",x"41"),
  2199 => (x"7f",x"7f",x"00",x"00"),
  2200 => (x"41",x"41",x"49",x"49"),
  2201 => (x"7f",x"7f",x"00",x"00"),
  2202 => (x"01",x"01",x"09",x"09"),
  2203 => (x"7f",x"3e",x"00",x"00"),
  2204 => (x"7a",x"7b",x"49",x"41"),
  2205 => (x"7f",x"7f",x"00",x"00"),
  2206 => (x"7f",x"7f",x"08",x"08"),
  2207 => (x"41",x"00",x"00",x"00"),
  2208 => (x"00",x"41",x"7f",x"7f"),
  2209 => (x"60",x"20",x"00",x"00"),
  2210 => (x"3f",x"7f",x"40",x"40"),
  2211 => (x"08",x"7f",x"7f",x"00"),
  2212 => (x"41",x"63",x"36",x"1c"),
  2213 => (x"7f",x"7f",x"00",x"00"),
  2214 => (x"40",x"40",x"40",x"40"),
  2215 => (x"06",x"7f",x"7f",x"00"),
  2216 => (x"7f",x"7f",x"06",x"0c"),
  2217 => (x"06",x"7f",x"7f",x"00"),
  2218 => (x"7f",x"7f",x"18",x"0c"),
  2219 => (x"7f",x"3e",x"00",x"00"),
  2220 => (x"3e",x"7f",x"41",x"41"),
  2221 => (x"7f",x"7f",x"00",x"00"),
  2222 => (x"06",x"0f",x"09",x"09"),
  2223 => (x"41",x"7f",x"3e",x"00"),
  2224 => (x"40",x"7e",x"7f",x"61"),
  2225 => (x"7f",x"7f",x"00",x"00"),
  2226 => (x"66",x"7f",x"19",x"09"),
  2227 => (x"6f",x"26",x"00",x"00"),
  2228 => (x"32",x"7b",x"59",x"4d"),
  2229 => (x"01",x"01",x"00",x"00"),
  2230 => (x"01",x"01",x"7f",x"7f"),
  2231 => (x"7f",x"3f",x"00",x"00"),
  2232 => (x"3f",x"7f",x"40",x"40"),
  2233 => (x"3f",x"0f",x"00",x"00"),
  2234 => (x"0f",x"3f",x"70",x"70"),
  2235 => (x"30",x"7f",x"7f",x"00"),
  2236 => (x"7f",x"7f",x"30",x"18"),
  2237 => (x"36",x"63",x"41",x"00"),
  2238 => (x"63",x"36",x"1c",x"1c"),
  2239 => (x"06",x"03",x"01",x"41"),
  2240 => (x"03",x"06",x"7c",x"7c"),
  2241 => (x"59",x"71",x"61",x"01"),
  2242 => (x"41",x"43",x"47",x"4d"),
  2243 => (x"7f",x"00",x"00",x"00"),
  2244 => (x"00",x"41",x"41",x"7f"),
  2245 => (x"06",x"03",x"01",x"00"),
  2246 => (x"60",x"30",x"18",x"0c"),
  2247 => (x"41",x"00",x"00",x"40"),
  2248 => (x"00",x"7f",x"7f",x"41"),
  2249 => (x"06",x"0c",x"08",x"00"),
  2250 => (x"08",x"0c",x"06",x"03"),
  2251 => (x"80",x"80",x"80",x"00"),
  2252 => (x"80",x"80",x"80",x"80"),
  2253 => (x"00",x"00",x"00",x"00"),
  2254 => (x"00",x"04",x"07",x"03"),
  2255 => (x"74",x"20",x"00",x"00"),
  2256 => (x"78",x"7c",x"54",x"54"),
  2257 => (x"7f",x"7f",x"00",x"00"),
  2258 => (x"38",x"7c",x"44",x"44"),
  2259 => (x"7c",x"38",x"00",x"00"),
  2260 => (x"00",x"44",x"44",x"44"),
  2261 => (x"7c",x"38",x"00",x"00"),
  2262 => (x"7f",x"7f",x"44",x"44"),
  2263 => (x"7c",x"38",x"00",x"00"),
  2264 => (x"18",x"5c",x"54",x"54"),
  2265 => (x"7e",x"04",x"00",x"00"),
  2266 => (x"00",x"05",x"05",x"7f"),
  2267 => (x"bc",x"18",x"00",x"00"),
  2268 => (x"7c",x"fc",x"a4",x"a4"),
  2269 => (x"7f",x"7f",x"00",x"00"),
  2270 => (x"78",x"7c",x"04",x"04"),
  2271 => (x"00",x"00",x"00",x"00"),
  2272 => (x"00",x"40",x"7d",x"3d"),
  2273 => (x"80",x"80",x"00",x"00"),
  2274 => (x"00",x"7d",x"fd",x"80"),
  2275 => (x"7f",x"7f",x"00",x"00"),
  2276 => (x"44",x"6c",x"38",x"10"),
  2277 => (x"00",x"00",x"00",x"00"),
  2278 => (x"00",x"40",x"7f",x"3f"),
  2279 => (x"0c",x"7c",x"7c",x"00"),
  2280 => (x"78",x"7c",x"0c",x"18"),
  2281 => (x"7c",x"7c",x"00",x"00"),
  2282 => (x"78",x"7c",x"04",x"04"),
  2283 => (x"7c",x"38",x"00",x"00"),
  2284 => (x"38",x"7c",x"44",x"44"),
  2285 => (x"fc",x"fc",x"00",x"00"),
  2286 => (x"18",x"3c",x"24",x"24"),
  2287 => (x"3c",x"18",x"00",x"00"),
  2288 => (x"fc",x"fc",x"24",x"24"),
  2289 => (x"7c",x"7c",x"00",x"00"),
  2290 => (x"08",x"0c",x"04",x"04"),
  2291 => (x"5c",x"48",x"00",x"00"),
  2292 => (x"20",x"74",x"54",x"54"),
  2293 => (x"3f",x"04",x"00",x"00"),
  2294 => (x"00",x"44",x"44",x"7f"),
  2295 => (x"7c",x"3c",x"00",x"00"),
  2296 => (x"7c",x"7c",x"40",x"40"),
  2297 => (x"3c",x"1c",x"00",x"00"),
  2298 => (x"1c",x"3c",x"60",x"60"),
  2299 => (x"60",x"7c",x"3c",x"00"),
  2300 => (x"3c",x"7c",x"60",x"30"),
  2301 => (x"38",x"6c",x"44",x"00"),
  2302 => (x"44",x"6c",x"38",x"10"),
  2303 => (x"bc",x"1c",x"00",x"00"),
  2304 => (x"1c",x"3c",x"60",x"e0"),
  2305 => (x"64",x"44",x"00",x"00"),
  2306 => (x"44",x"4c",x"5c",x"74"),
  2307 => (x"08",x"08",x"00",x"00"),
  2308 => (x"41",x"41",x"77",x"3e"),
  2309 => (x"00",x"00",x"00",x"00"),
  2310 => (x"00",x"00",x"7f",x"7f"),
  2311 => (x"41",x"41",x"00",x"00"),
  2312 => (x"08",x"08",x"3e",x"77"),
  2313 => (x"01",x"01",x"02",x"00"),
  2314 => (x"01",x"02",x"02",x"03"),
  2315 => (x"7f",x"7f",x"7f",x"00"),
  2316 => (x"7f",x"7f",x"7f",x"7f"),
  2317 => (x"1c",x"08",x"08",x"00"),
  2318 => (x"7f",x"3e",x"3e",x"1c"),
  2319 => (x"3e",x"7f",x"7f",x"7f"),
  2320 => (x"08",x"1c",x"1c",x"3e"),
  2321 => (x"18",x"10",x"00",x"08"),
  2322 => (x"10",x"18",x"7c",x"7c"),
  2323 => (x"30",x"10",x"00",x"00"),
  2324 => (x"10",x"30",x"7c",x"7c"),
  2325 => (x"60",x"30",x"10",x"00"),
  2326 => (x"06",x"1e",x"78",x"60"),
  2327 => (x"3c",x"66",x"42",x"00"),
  2328 => (x"42",x"66",x"3c",x"18"),
  2329 => (x"6a",x"38",x"78",x"00"),
  2330 => (x"38",x"6c",x"c6",x"c2"),
  2331 => (x"00",x"00",x"60",x"00"),
  2332 => (x"60",x"00",x"00",x"60"),
  2333 => (x"5b",x"5e",x"0e",x"00"),
  2334 => (x"1e",x"0e",x"5d",x"5c"),
  2335 => (x"fa",x"c2",x"4c",x"71"),
  2336 => (x"c0",x"4d",x"bf",x"c1"),
  2337 => (x"74",x"1e",x"c0",x"4b"),
  2338 => (x"87",x"c7",x"02",x"ab"),
  2339 => (x"c0",x"48",x"a6",x"c4"),
  2340 => (x"c4",x"87",x"c5",x"78"),
  2341 => (x"78",x"c1",x"48",x"a6"),
  2342 => (x"73",x"1e",x"66",x"c4"),
  2343 => (x"87",x"df",x"ee",x"49"),
  2344 => (x"e0",x"c0",x"86",x"c8"),
  2345 => (x"87",x"ef",x"ef",x"49"),
  2346 => (x"6a",x"4a",x"a5",x"c4"),
  2347 => (x"87",x"f0",x"f0",x"49"),
  2348 => (x"cb",x"87",x"c6",x"f1"),
  2349 => (x"c8",x"83",x"c1",x"85"),
  2350 => (x"ff",x"04",x"ab",x"b7"),
  2351 => (x"26",x"26",x"87",x"c7"),
  2352 => (x"26",x"4c",x"26",x"4d"),
  2353 => (x"1e",x"4f",x"26",x"4b"),
  2354 => (x"fa",x"c2",x"4a",x"71"),
  2355 => (x"fa",x"c2",x"5a",x"c5"),
  2356 => (x"78",x"c7",x"48",x"c5"),
  2357 => (x"87",x"dd",x"fe",x"49"),
  2358 => (x"73",x"1e",x"4f",x"26"),
  2359 => (x"c0",x"4a",x"71",x"1e"),
  2360 => (x"d3",x"03",x"aa",x"b7"),
  2361 => (x"fa",x"e0",x"c2",x"87"),
  2362 => (x"87",x"c4",x"05",x"bf"),
  2363 => (x"87",x"c2",x"4b",x"c1"),
  2364 => (x"e0",x"c2",x"4b",x"c0"),
  2365 => (x"87",x"c4",x"5b",x"fe"),
  2366 => (x"5a",x"fe",x"e0",x"c2"),
  2367 => (x"bf",x"fa",x"e0",x"c2"),
  2368 => (x"c1",x"9a",x"c1",x"4a"),
  2369 => (x"ec",x"49",x"a2",x"c0"),
  2370 => (x"48",x"fc",x"87",x"e8"),
  2371 => (x"bf",x"fa",x"e0",x"c2"),
  2372 => (x"87",x"ef",x"fe",x"78"),
  2373 => (x"c4",x"4a",x"71",x"1e"),
  2374 => (x"49",x"72",x"1e",x"66"),
  2375 => (x"87",x"dd",x"df",x"ff"),
  2376 => (x"1e",x"4f",x"26",x"26"),
  2377 => (x"bf",x"fa",x"e0",x"c2"),
  2378 => (x"cd",x"dc",x"ff",x"49"),
  2379 => (x"f9",x"f9",x"c2",x"87"),
  2380 => (x"78",x"bf",x"e8",x"48"),
  2381 => (x"48",x"f5",x"f9",x"c2"),
  2382 => (x"c2",x"78",x"bf",x"ec"),
  2383 => (x"4a",x"bf",x"f9",x"f9"),
  2384 => (x"99",x"ff",x"c3",x"49"),
  2385 => (x"72",x"2a",x"b7",x"c8"),
  2386 => (x"c2",x"b0",x"71",x"48"),
  2387 => (x"26",x"58",x"c1",x"fa"),
  2388 => (x"5b",x"5e",x"0e",x"4f"),
  2389 => (x"71",x"0e",x"5d",x"5c"),
  2390 => (x"87",x"c7",x"ff",x"4b"),
  2391 => (x"48",x"f4",x"f9",x"c2"),
  2392 => (x"49",x"73",x"50",x"c0"),
  2393 => (x"87",x"f2",x"db",x"ff"),
  2394 => (x"c2",x"4c",x"49",x"70"),
  2395 => (x"49",x"ee",x"cb",x"9c"),
  2396 => (x"70",x"87",x"cf",x"cb"),
  2397 => (x"f9",x"c2",x"4d",x"49"),
  2398 => (x"05",x"bf",x"97",x"f4"),
  2399 => (x"d0",x"87",x"e4",x"c1"),
  2400 => (x"f9",x"c2",x"49",x"66"),
  2401 => (x"05",x"99",x"bf",x"fd"),
  2402 => (x"66",x"d4",x"87",x"d7"),
  2403 => (x"f5",x"f9",x"c2",x"49"),
  2404 => (x"cc",x"05",x"99",x"bf"),
  2405 => (x"ff",x"49",x"73",x"87"),
  2406 => (x"70",x"87",x"ff",x"da"),
  2407 => (x"c2",x"c1",x"02",x"98"),
  2408 => (x"fd",x"4c",x"c1",x"87"),
  2409 => (x"49",x"75",x"87",x"fd"),
  2410 => (x"70",x"87",x"e3",x"ca"),
  2411 => (x"87",x"c6",x"02",x"98"),
  2412 => (x"48",x"f4",x"f9",x"c2"),
  2413 => (x"f9",x"c2",x"50",x"c1"),
  2414 => (x"05",x"bf",x"97",x"f4"),
  2415 => (x"c2",x"87",x"e4",x"c0"),
  2416 => (x"49",x"bf",x"fd",x"f9"),
  2417 => (x"05",x"99",x"66",x"d0"),
  2418 => (x"c2",x"87",x"d6",x"ff"),
  2419 => (x"49",x"bf",x"f5",x"f9"),
  2420 => (x"05",x"99",x"66",x"d4"),
  2421 => (x"73",x"87",x"ca",x"ff"),
  2422 => (x"fd",x"d9",x"ff",x"49"),
  2423 => (x"05",x"98",x"70",x"87"),
  2424 => (x"74",x"87",x"fe",x"fe"),
  2425 => (x"87",x"d7",x"fb",x"48"),
  2426 => (x"5c",x"5b",x"5e",x"0e"),
  2427 => (x"86",x"f4",x"0e",x"5d"),
  2428 => (x"ec",x"4c",x"4d",x"c0"),
  2429 => (x"a6",x"c4",x"7e",x"bf"),
  2430 => (x"c1",x"fa",x"c2",x"48"),
  2431 => (x"1e",x"c1",x"78",x"bf"),
  2432 => (x"49",x"c7",x"1e",x"c0"),
  2433 => (x"c8",x"87",x"ca",x"fd"),
  2434 => (x"02",x"98",x"70",x"86"),
  2435 => (x"49",x"ff",x"87",x"ce"),
  2436 => (x"c1",x"87",x"c7",x"fb"),
  2437 => (x"d9",x"ff",x"49",x"da"),
  2438 => (x"4d",x"c1",x"87",x"c0"),
  2439 => (x"97",x"f4",x"f9",x"c2"),
  2440 => (x"87",x"c3",x"02",x"bf"),
  2441 => (x"c2",x"87",x"c0",x"c9"),
  2442 => (x"4b",x"bf",x"f9",x"f9"),
  2443 => (x"bf",x"fa",x"e0",x"c2"),
  2444 => (x"87",x"eb",x"c0",x"05"),
  2445 => (x"ff",x"49",x"fd",x"c3"),
  2446 => (x"c3",x"87",x"df",x"d8"),
  2447 => (x"d8",x"ff",x"49",x"fa"),
  2448 => (x"49",x"73",x"87",x"d8"),
  2449 => (x"71",x"99",x"ff",x"c3"),
  2450 => (x"fb",x"49",x"c0",x"1e"),
  2451 => (x"49",x"73",x"87",x"c6"),
  2452 => (x"71",x"29",x"b7",x"c8"),
  2453 => (x"fa",x"49",x"c1",x"1e"),
  2454 => (x"86",x"c8",x"87",x"fa"),
  2455 => (x"c2",x"87",x"c1",x"c6"),
  2456 => (x"4b",x"bf",x"fd",x"f9"),
  2457 => (x"87",x"dd",x"02",x"9b"),
  2458 => (x"bf",x"f6",x"e0",x"c2"),
  2459 => (x"87",x"de",x"c7",x"49"),
  2460 => (x"c4",x"05",x"98",x"70"),
  2461 => (x"d2",x"4b",x"c0",x"87"),
  2462 => (x"49",x"e0",x"c2",x"87"),
  2463 => (x"c2",x"87",x"c3",x"c7"),
  2464 => (x"c6",x"58",x"fa",x"e0"),
  2465 => (x"f6",x"e0",x"c2",x"87"),
  2466 => (x"73",x"78",x"c0",x"48"),
  2467 => (x"05",x"99",x"c2",x"49"),
  2468 => (x"eb",x"c3",x"87",x"ce"),
  2469 => (x"c1",x"d7",x"ff",x"49"),
  2470 => (x"c2",x"49",x"70",x"87"),
  2471 => (x"87",x"c2",x"02",x"99"),
  2472 => (x"49",x"73",x"4c",x"fb"),
  2473 => (x"ce",x"05",x"99",x"c1"),
  2474 => (x"49",x"f4",x"c3",x"87"),
  2475 => (x"87",x"ea",x"d6",x"ff"),
  2476 => (x"99",x"c2",x"49",x"70"),
  2477 => (x"fa",x"87",x"c2",x"02"),
  2478 => (x"c8",x"49",x"73",x"4c"),
  2479 => (x"87",x"ce",x"05",x"99"),
  2480 => (x"ff",x"49",x"f5",x"c3"),
  2481 => (x"70",x"87",x"d3",x"d6"),
  2482 => (x"02",x"99",x"c2",x"49"),
  2483 => (x"fa",x"c2",x"87",x"d5"),
  2484 => (x"ca",x"02",x"bf",x"c5"),
  2485 => (x"88",x"c1",x"48",x"87"),
  2486 => (x"58",x"c9",x"fa",x"c2"),
  2487 => (x"ff",x"87",x"c2",x"c0"),
  2488 => (x"73",x"4d",x"c1",x"4c"),
  2489 => (x"05",x"99",x"c4",x"49"),
  2490 => (x"f2",x"c3",x"87",x"ce"),
  2491 => (x"e9",x"d5",x"ff",x"49"),
  2492 => (x"c2",x"49",x"70",x"87"),
  2493 => (x"87",x"dc",x"02",x"99"),
  2494 => (x"bf",x"c5",x"fa",x"c2"),
  2495 => (x"b7",x"c7",x"48",x"7e"),
  2496 => (x"cb",x"c0",x"03",x"a8"),
  2497 => (x"c1",x"48",x"6e",x"87"),
  2498 => (x"c9",x"fa",x"c2",x"80"),
  2499 => (x"87",x"c2",x"c0",x"58"),
  2500 => (x"4d",x"c1",x"4c",x"fe"),
  2501 => (x"ff",x"49",x"fd",x"c3"),
  2502 => (x"70",x"87",x"ff",x"d4"),
  2503 => (x"02",x"99",x"c2",x"49"),
  2504 => (x"c2",x"87",x"d5",x"c0"),
  2505 => (x"02",x"bf",x"c5",x"fa"),
  2506 => (x"c2",x"87",x"c9",x"c0"),
  2507 => (x"c0",x"48",x"c5",x"fa"),
  2508 => (x"87",x"c2",x"c0",x"78"),
  2509 => (x"4d",x"c1",x"4c",x"fd"),
  2510 => (x"ff",x"49",x"fa",x"c3"),
  2511 => (x"70",x"87",x"db",x"d4"),
  2512 => (x"02",x"99",x"c2",x"49"),
  2513 => (x"c2",x"87",x"d9",x"c0"),
  2514 => (x"48",x"bf",x"c5",x"fa"),
  2515 => (x"03",x"a8",x"b7",x"c7"),
  2516 => (x"c2",x"87",x"c9",x"c0"),
  2517 => (x"c7",x"48",x"c5",x"fa"),
  2518 => (x"87",x"c2",x"c0",x"78"),
  2519 => (x"4d",x"c1",x"4c",x"fc"),
  2520 => (x"03",x"ac",x"b7",x"c0"),
  2521 => (x"c4",x"87",x"d1",x"c0"),
  2522 => (x"d8",x"c1",x"4a",x"66"),
  2523 => (x"c0",x"02",x"6a",x"82"),
  2524 => (x"4b",x"6a",x"87",x"c6"),
  2525 => (x"0f",x"73",x"49",x"74"),
  2526 => (x"f0",x"c3",x"1e",x"c0"),
  2527 => (x"49",x"da",x"c1",x"1e"),
  2528 => (x"c8",x"87",x"ce",x"f7"),
  2529 => (x"02",x"98",x"70",x"86"),
  2530 => (x"c8",x"87",x"e2",x"c0"),
  2531 => (x"fa",x"c2",x"48",x"a6"),
  2532 => (x"c8",x"78",x"bf",x"c5"),
  2533 => (x"91",x"cb",x"49",x"66"),
  2534 => (x"71",x"48",x"66",x"c4"),
  2535 => (x"6e",x"7e",x"70",x"80"),
  2536 => (x"c8",x"c0",x"02",x"bf"),
  2537 => (x"4b",x"bf",x"6e",x"87"),
  2538 => (x"73",x"49",x"66",x"c8"),
  2539 => (x"02",x"9d",x"75",x"0f"),
  2540 => (x"c2",x"87",x"c8",x"c0"),
  2541 => (x"49",x"bf",x"c5",x"fa"),
  2542 => (x"c2",x"87",x"fa",x"f2"),
  2543 => (x"02",x"bf",x"fe",x"e0"),
  2544 => (x"49",x"87",x"dd",x"c0"),
  2545 => (x"70",x"87",x"c7",x"c2"),
  2546 => (x"d3",x"c0",x"02",x"98"),
  2547 => (x"c5",x"fa",x"c2",x"87"),
  2548 => (x"e0",x"f2",x"49",x"bf"),
  2549 => (x"f4",x"49",x"c0",x"87"),
  2550 => (x"e0",x"c2",x"87",x"c0"),
  2551 => (x"78",x"c0",x"48",x"fe"),
  2552 => (x"da",x"f3",x"8e",x"f4"),
  2553 => (x"5b",x"5e",x"0e",x"87"),
  2554 => (x"1e",x"0e",x"5d",x"5c"),
  2555 => (x"fa",x"c2",x"4c",x"71"),
  2556 => (x"c1",x"49",x"bf",x"c1"),
  2557 => (x"c1",x"4d",x"a1",x"cd"),
  2558 => (x"7e",x"69",x"81",x"d1"),
  2559 => (x"cf",x"02",x"9c",x"74"),
  2560 => (x"4b",x"a5",x"c4",x"87"),
  2561 => (x"fa",x"c2",x"7b",x"74"),
  2562 => (x"f2",x"49",x"bf",x"c1"),
  2563 => (x"7b",x"6e",x"87",x"f9"),
  2564 => (x"c4",x"05",x"9c",x"74"),
  2565 => (x"c2",x"4b",x"c0",x"87"),
  2566 => (x"73",x"4b",x"c1",x"87"),
  2567 => (x"87",x"fa",x"f2",x"49"),
  2568 => (x"c7",x"02",x"66",x"d4"),
  2569 => (x"87",x"da",x"49",x"87"),
  2570 => (x"87",x"c2",x"4a",x"70"),
  2571 => (x"e1",x"c2",x"4a",x"c0"),
  2572 => (x"f2",x"26",x"5a",x"c2"),
  2573 => (x"00",x"00",x"87",x"c9"),
  2574 => (x"00",x"00",x"00",x"00"),
  2575 => (x"00",x"00",x"00",x"00"),
  2576 => (x"71",x"1e",x"00",x"00"),
  2577 => (x"bf",x"c8",x"ff",x"4a"),
  2578 => (x"48",x"a1",x"72",x"49"),
  2579 => (x"ff",x"1e",x"4f",x"26"),
  2580 => (x"fe",x"89",x"bf",x"c8"),
  2581 => (x"c0",x"c0",x"c0",x"c0"),
  2582 => (x"c4",x"01",x"a9",x"c0"),
  2583 => (x"c2",x"4a",x"c0",x"87"),
  2584 => (x"72",x"4a",x"c1",x"87"),
  2585 => (x"1e",x"4f",x"26",x"48"),
  2586 => (x"bf",x"f5",x"e2",x"c2"),
  2587 => (x"c2",x"b9",x"c1",x"49"),
  2588 => (x"ff",x"59",x"f9",x"e2"),
  2589 => (x"ff",x"c3",x"48",x"d4"),
  2590 => (x"48",x"d0",x"ff",x"78"),
  2591 => (x"ff",x"78",x"e1",x"c0"),
  2592 => (x"78",x"c1",x"48",x"d4"),
  2593 => (x"78",x"71",x"31",x"c4"),
  2594 => (x"c0",x"48",x"d0",x"ff"),
  2595 => (x"4f",x"26",x"78",x"e0"),
  2596 => (x"e9",x"e2",x"c2",x"1e"),
  2597 => (x"e8",x"f4",x"c2",x"1e"),
  2598 => (x"d4",x"fd",x"fd",x"49"),
  2599 => (x"70",x"86",x"c4",x"87"),
  2600 => (x"87",x"c3",x"02",x"98"),
  2601 => (x"26",x"87",x"c0",x"ff"),
  2602 => (x"4b",x"35",x"31",x"4f"),
  2603 => (x"20",x"20",x"5a",x"48"),
  2604 => (x"47",x"46",x"43",x"20"),
  2605 => (x"00",x"00",x"00",x"00"),
  2606 => (x"5b",x"5e",x"0e",x"00"),
  2607 => (x"c2",x"0e",x"5d",x"5c"),
  2608 => (x"4a",x"bf",x"f5",x"f9"),
  2609 => (x"bf",x"e2",x"e4",x"c2"),
  2610 => (x"bc",x"72",x"4c",x"49"),
  2611 => (x"c6",x"ff",x"4d",x"71"),
  2612 => (x"4b",x"c0",x"87",x"de"),
  2613 => (x"99",x"d0",x"49",x"74"),
  2614 => (x"87",x"e7",x"c0",x"02"),
  2615 => (x"c8",x"48",x"d0",x"ff"),
  2616 => (x"d4",x"ff",x"78",x"e1"),
  2617 => (x"75",x"78",x"c5",x"48"),
  2618 => (x"02",x"99",x"d0",x"49"),
  2619 => (x"f0",x"c3",x"87",x"c3"),
  2620 => (x"c3",x"e7",x"c2",x"78"),
  2621 => (x"11",x"81",x"73",x"49"),
  2622 => (x"08",x"d4",x"ff",x"48"),
  2623 => (x"48",x"d0",x"ff",x"78"),
  2624 => (x"c1",x"78",x"e0",x"c0"),
  2625 => (x"c8",x"83",x"2d",x"2c"),
  2626 => (x"c7",x"ff",x"04",x"ab"),
  2627 => (x"d7",x"c5",x"ff",x"87"),
  2628 => (x"e2",x"e4",x"c2",x"87"),
  2629 => (x"f5",x"f9",x"c2",x"48"),
  2630 => (x"4d",x"26",x"78",x"bf"),
  2631 => (x"4b",x"26",x"4c",x"26"),
  2632 => (x"00",x"00",x"4f",x"26"),
  2633 => (x"c1",x"1e",x"00",x"00"),
  2634 => (x"de",x"48",x"d7",x"e7"),
  2635 => (x"c2",x"1e",x"c8",x"50"),
  2636 => (x"fe",x"49",x"c9",x"fa"),
  2637 => (x"c4",x"87",x"c5",x"d5"),
  2638 => (x"c2",x"1e",x"72",x"86"),
  2639 => (x"c2",x"48",x"cc",x"e6"),
  2640 => (x"c4",x"49",x"d1",x"fa"),
  2641 => (x"41",x"20",x"4a",x"a1"),
  2642 => (x"f9",x"05",x"aa",x"71"),
  2643 => (x"c2",x"4a",x"26",x"87"),
  2644 => (x"fd",x"49",x"d0",x"e6"),
  2645 => (x"70",x"87",x"fb",x"f8"),
  2646 => (x"c5",x"02",x"9a",x"4a"),
  2647 => (x"c7",x"fe",x"49",x"87"),
  2648 => (x"1e",x"72",x"87",x"e4"),
  2649 => (x"48",x"dc",x"e6",x"c2"),
  2650 => (x"49",x"d1",x"fa",x"c2"),
  2651 => (x"20",x"4a",x"a1",x"c4"),
  2652 => (x"05",x"aa",x"71",x"41"),
  2653 => (x"4a",x"26",x"87",x"f9"),
  2654 => (x"49",x"c9",x"fa",x"c2"),
  2655 => (x"87",x"d5",x"d9",x"fe"),
  2656 => (x"c5",x"fe",x"49",x"c0"),
  2657 => (x"e6",x"c2",x"87",x"e2"),
  2658 => (x"4f",x"26",x"48",x"e0"),
  2659 => (x"00",x"20",x"20",x"20"),
  2660 => (x"45",x"54",x"4f",x"4a"),
  2661 => (x"20",x"20",x"4f",x"47"),
  2662 => (x"00",x"20",x"20",x"20"),
  2663 => (x"00",x"43",x"52",x"41"),
  2664 => (x"20",x"43",x"52",x"41"),
  2665 => (x"20",x"74",x"6f",x"6e"),
  2666 => (x"6e",x"75",x"6f",x"66"),
  2667 => (x"4c",x"20",x"2e",x"64"),
  2668 => (x"20",x"64",x"61",x"6f"),
  2669 => (x"00",x"43",x"52",x"41"),
  2670 => (x"87",x"ec",x"f0",x"1e"),
  2671 => (x"f8",x"87",x"fa",x"fb"),
  2672 => (x"16",x"4f",x"26",x"87"),
  2673 => (x"2e",x"25",x"26",x"1e"),
  2674 => (x"2e",x"3e",x"3d",x"36"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

